library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"78e0c048",
     1 => x"1e4f2626",
     2 => x"b7c24a71",
     3 => x"87c303aa",
     4 => x"ce87c282",
     5 => x"1e66c482",
     6 => x"d5ff4972",
     7 => x"4f262687",
     8 => x"4ad4ff1e",
     9 => x"ff7affc3",
    10 => x"e1c848d0",
    11 => x"c37ade78",
    12 => x"7abfd3c5",
    13 => x"28c84849",
    14 => x"48717a70",
    15 => x"7a7028d0",
    16 => x"28d84871",
    17 => x"c5c37a70",
    18 => x"497abfd7",
    19 => x"7028c848",
    20 => x"d048717a",
    21 => x"717a7028",
    22 => x"7028d848",
    23 => x"48d0ff7a",
    24 => x"2678e0c0",
    25 => x"1e731e4f",
    26 => x"c5c34a71",
    27 => x"724bbfd3",
    28 => x"aae0c02b",
    29 => x"7287ce04",
    30 => x"89e0c049",
    31 => x"bfd7c5c3",
    32 => x"cf2b714b",
    33 => x"49e0c087",
    34 => x"c5c38972",
    35 => x"7148bfd7",
    36 => x"b3497030",
    37 => x"739b66c8",
    38 => x"2687c448",
    39 => x"264c264d",
    40 => x"0e4f264b",
    41 => x"5d5c5b5e",
    42 => x"7186ec0e",
    43 => x"d3c5c34b",
    44 => x"734c7ebf",
    45 => x"abe0c02c",
    46 => x"87e0c004",
    47 => x"c048a6c4",
    48 => x"c0497378",
    49 => x"4a7189e0",
    50 => x"4866e4c0",
    51 => x"a6cc3072",
    52 => x"d7c5c358",
    53 => x"714c4dbf",
    54 => x"87e4c02c",
    55 => x"e4c04973",
    56 => x"30714866",
    57 => x"c058a6c8",
    58 => x"897349e0",
    59 => x"4866e4c0",
    60 => x"a6cc2871",
    61 => x"d7c5c358",
    62 => x"71484dbf",
    63 => x"b4497030",
    64 => x"9c66e4c0",
    65 => x"e8c084c1",
    66 => x"c204ac66",
    67 => x"c04cc087",
    68 => x"d304abe0",
    69 => x"48a6cc87",
    70 => x"497378c0",
    71 => x"7489e0c0",
    72 => x"d4307148",
    73 => x"87d558a6",
    74 => x"48744973",
    75 => x"a6d03071",
    76 => x"49e0c058",
    77 => x"48748973",
    78 => x"a6d42871",
    79 => x"4a66c458",
    80 => x"9a6ebaff",
    81 => x"ff4966c8",
    82 => x"729975b9",
    83 => x"b066cc48",
    84 => x"58d7c5c3",
    85 => x"66d04871",
    86 => x"dbc5c3b0",
    87 => x"87c0fb58",
    88 => x"f6fc8eec",
    89 => x"d0ff1e87",
    90 => x"78c9c848",
    91 => x"d4ff4871",
    92 => x"4f267808",
    93 => x"494a711e",
    94 => x"d0ff87eb",
    95 => x"2678c848",
    96 => x"1e731e4f",
    97 => x"c5c34b71",
    98 => x"c302bfe7",
    99 => x"87ebc287",
   100 => x"c848d0ff",
   101 => x"497378c9",
   102 => x"ffb1e0c0",
   103 => x"787148d4",
   104 => x"48dbc5c3",
   105 => x"66c878c0",
   106 => x"c387c502",
   107 => x"87c249ff",
   108 => x"c5c349c0",
   109 => x"66cc59e3",
   110 => x"c587c602",
   111 => x"c44ad5d5",
   112 => x"ffffcf87",
   113 => x"e7c5c34a",
   114 => x"e7c5c35a",
   115 => x"c478c148",
   116 => x"264d2687",
   117 => x"264b264c",
   118 => x"5b5e0e4f",
   119 => x"710e5d5c",
   120 => x"e3c5c34a",
   121 => x"9a724cbf",
   122 => x"4987cb02",
   123 => x"c5c291c8",
   124 => x"83714bf7",
   125 => x"c9c287c4",
   126 => x"4dc04bf7",
   127 => x"99744913",
   128 => x"bfdfc5c3",
   129 => x"48d4ffb9",
   130 => x"b7c17871",
   131 => x"b7c8852c",
   132 => x"87e804ad",
   133 => x"bfdbc5c3",
   134 => x"c380c848",
   135 => x"fe58dfc5",
   136 => x"731e87ef",
   137 => x"134b711e",
   138 => x"cb029a4a",
   139 => x"fe497287",
   140 => x"4a1387e7",
   141 => x"87f5059a",
   142 => x"1e87dafe",
   143 => x"bfdbc5c3",
   144 => x"dbc5c349",
   145 => x"78a1c148",
   146 => x"a9b7c0c4",
   147 => x"ff87db03",
   148 => x"c5c348d4",
   149 => x"c378bfdf",
   150 => x"49bfdbc5",
   151 => x"48dbc5c3",
   152 => x"c478a1c1",
   153 => x"04a9b7c0",
   154 => x"d0ff87e5",
   155 => x"c378c848",
   156 => x"c048e7c5",
   157 => x"004f2678",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"5f5f0000",
   161 => x"00000000",
   162 => x"03000303",
   163 => x"14000003",
   164 => x"7f147f7f",
   165 => x"0000147f",
   166 => x"6b6b2e24",
   167 => x"4c00123a",
   168 => x"6c18366a",
   169 => x"30003256",
   170 => x"77594f7e",
   171 => x"0040683a",
   172 => x"03070400",
   173 => x"00000000",
   174 => x"633e1c00",
   175 => x"00000041",
   176 => x"3e634100",
   177 => x"0800001c",
   178 => x"1c1c3e2a",
   179 => x"00082a3e",
   180 => x"3e3e0808",
   181 => x"00000808",
   182 => x"60e08000",
   183 => x"00000000",
   184 => x"08080808",
   185 => x"00000808",
   186 => x"60600000",
   187 => x"40000000",
   188 => x"0c183060",
   189 => x"00010306",
   190 => x"4d597f3e",
   191 => x"00003e7f",
   192 => x"7f7f0604",
   193 => x"00000000",
   194 => x"59716342",
   195 => x"0000464f",
   196 => x"49496322",
   197 => x"1800367f",
   198 => x"7f13161c",
   199 => x"0000107f",
   200 => x"45456727",
   201 => x"0000397d",
   202 => x"494b7e3c",
   203 => x"00003079",
   204 => x"79710101",
   205 => x"0000070f",
   206 => x"49497f36",
   207 => x"0000367f",
   208 => x"69494f06",
   209 => x"00001e3f",
   210 => x"66660000",
   211 => x"00000000",
   212 => x"66e68000",
   213 => x"00000000",
   214 => x"14140808",
   215 => x"00002222",
   216 => x"14141414",
   217 => x"00001414",
   218 => x"14142222",
   219 => x"00000808",
   220 => x"59510302",
   221 => x"3e00060f",
   222 => x"555d417f",
   223 => x"00001e1f",
   224 => x"09097f7e",
   225 => x"00007e7f",
   226 => x"49497f7f",
   227 => x"0000367f",
   228 => x"41633e1c",
   229 => x"00004141",
   230 => x"63417f7f",
   231 => x"00001c3e",
   232 => x"49497f7f",
   233 => x"00004141",
   234 => x"09097f7f",
   235 => x"00000101",
   236 => x"49417f3e",
   237 => x"00007a7b",
   238 => x"08087f7f",
   239 => x"00007f7f",
   240 => x"7f7f4100",
   241 => x"00000041",
   242 => x"40406020",
   243 => x"7f003f7f",
   244 => x"361c087f",
   245 => x"00004163",
   246 => x"40407f7f",
   247 => x"7f004040",
   248 => x"060c067f",
   249 => x"7f007f7f",
   250 => x"180c067f",
   251 => x"00007f7f",
   252 => x"41417f3e",
   253 => x"00003e7f",
   254 => x"09097f7f",
   255 => x"3e00060f",
   256 => x"7f61417f",
   257 => x"0000407e",
   258 => x"19097f7f",
   259 => x"0000667f",
   260 => x"594d6f26",
   261 => x"0000327b",
   262 => x"7f7f0101",
   263 => x"00000101",
   264 => x"40407f3f",
   265 => x"00003f7f",
   266 => x"70703f0f",
   267 => x"7f000f3f",
   268 => x"3018307f",
   269 => x"41007f7f",
   270 => x"1c1c3663",
   271 => x"01416336",
   272 => x"7c7c0603",
   273 => x"61010306",
   274 => x"474d5971",
   275 => x"00004143",
   276 => x"417f7f00",
   277 => x"01000041",
   278 => x"180c0603",
   279 => x"00406030",
   280 => x"7f414100",
   281 => x"0800007f",
   282 => x"0603060c",
   283 => x"8000080c",
   284 => x"80808080",
   285 => x"00008080",
   286 => x"07030000",
   287 => x"00000004",
   288 => x"54547420",
   289 => x"0000787c",
   290 => x"44447f7f",
   291 => x"0000387c",
   292 => x"44447c38",
   293 => x"00000044",
   294 => x"44447c38",
   295 => x"00007f7f",
   296 => x"54547c38",
   297 => x"0000185c",
   298 => x"057f7e04",
   299 => x"00000005",
   300 => x"a4a4bc18",
   301 => x"00007cfc",
   302 => x"04047f7f",
   303 => x"0000787c",
   304 => x"7d3d0000",
   305 => x"00000040",
   306 => x"fd808080",
   307 => x"0000007d",
   308 => x"38107f7f",
   309 => x"0000446c",
   310 => x"7f3f0000",
   311 => x"7c000040",
   312 => x"0c180c7c",
   313 => x"0000787c",
   314 => x"04047c7c",
   315 => x"0000787c",
   316 => x"44447c38",
   317 => x"0000387c",
   318 => x"2424fcfc",
   319 => x"0000183c",
   320 => x"24243c18",
   321 => x"0000fcfc",
   322 => x"04047c7c",
   323 => x"0000080c",
   324 => x"54545c48",
   325 => x"00002074",
   326 => x"447f3f04",
   327 => x"00000044",
   328 => x"40407c3c",
   329 => x"00007c7c",
   330 => x"60603c1c",
   331 => x"3c001c3c",
   332 => x"6030607c",
   333 => x"44003c7c",
   334 => x"3810386c",
   335 => x"0000446c",
   336 => x"60e0bc1c",
   337 => x"00001c3c",
   338 => x"5c746444",
   339 => x"0000444c",
   340 => x"773e0808",
   341 => x"00004141",
   342 => x"7f7f0000",
   343 => x"00000000",
   344 => x"3e774141",
   345 => x"02000808",
   346 => x"02030101",
   347 => x"7f000102",
   348 => x"7f7f7f7f",
   349 => x"08007f7f",
   350 => x"3e1c1c08",
   351 => x"7f7f7f3e",
   352 => x"1c3e3e7f",
   353 => x"0008081c",
   354 => x"7c7c1810",
   355 => x"00001018",
   356 => x"7c7c3010",
   357 => x"10001030",
   358 => x"78606030",
   359 => x"4200061e",
   360 => x"3c183c66",
   361 => x"78004266",
   362 => x"c6c26a38",
   363 => x"6000386c",
   364 => x"00600000",
   365 => x"0e006000",
   366 => x"5d5c5b5e",
   367 => x"4c711e0e",
   368 => x"bff8c5c3",
   369 => x"c04bc04d",
   370 => x"02ab741e",
   371 => x"a6c487c7",
   372 => x"c578c048",
   373 => x"48a6c487",
   374 => x"66c478c1",
   375 => x"ee49731e",
   376 => x"86c887df",
   377 => x"ef49e0c0",
   378 => x"a5c487ef",
   379 => x"f0496a4a",
   380 => x"c6f187f0",
   381 => x"c185cb87",
   382 => x"abb7c883",
   383 => x"87c7ff04",
   384 => x"264d2626",
   385 => x"264b264c",
   386 => x"4a711e4f",
   387 => x"5afcc5c3",
   388 => x"48fcc5c3",
   389 => x"fe4978c7",
   390 => x"4f2687dd",
   391 => x"711e731e",
   392 => x"aab7c04a",
   393 => x"c287d303",
   394 => x"05bffbe5",
   395 => x"4bc187c4",
   396 => x"4bc087c2",
   397 => x"5bffe5c2",
   398 => x"e5c287c4",
   399 => x"e5c25aff",
   400 => x"c14abffb",
   401 => x"a2c0c19a",
   402 => x"87e8ec49",
   403 => x"e5c248fc",
   404 => x"fe78bffb",
   405 => x"711e87ef",
   406 => x"1e66c44a",
   407 => x"e6e64972",
   408 => x"4f262687",
   409 => x"fbe5c21e",
   410 => x"daff49bf",
   411 => x"c5c387f6",
   412 => x"bfe848f0",
   413 => x"ecc5c378",
   414 => x"78bfec48",
   415 => x"bff0c5c3",
   416 => x"ffc3494a",
   417 => x"2ab7c899",
   418 => x"b0714872",
   419 => x"58f8c5c3",
   420 => x"5e0e4f26",
   421 => x"0e5d5c5b",
   422 => x"c7ff4b71",
   423 => x"ebc5c387",
   424 => x"7350c048",
   425 => x"dbdaff49",
   426 => x"4c497087",
   427 => x"eecb9cc2",
   428 => x"87cfcb49",
   429 => x"c34d4970",
   430 => x"bf97ebc5",
   431 => x"87e4c105",
   432 => x"c34966d0",
   433 => x"99bff4c5",
   434 => x"d487d705",
   435 => x"c5c34966",
   436 => x"0599bfec",
   437 => x"497387cc",
   438 => x"87e8d9ff",
   439 => x"c1029870",
   440 => x"4cc187c2",
   441 => x"7587fdfd",
   442 => x"87e3ca49",
   443 => x"c6029870",
   444 => x"ebc5c387",
   445 => x"c350c148",
   446 => x"bf97ebc5",
   447 => x"87e4c005",
   448 => x"bff4c5c3",
   449 => x"9966d049",
   450 => x"87d6ff05",
   451 => x"bfecc5c3",
   452 => x"9966d449",
   453 => x"87caff05",
   454 => x"d8ff4973",
   455 => x"987087e6",
   456 => x"87fefe05",
   457 => x"d8fb4874",
   458 => x"5b5e0e87",
   459 => x"f40e5d5c",
   460 => x"4c4dc086",
   461 => x"c47ebfec",
   462 => x"c5c348a6",
   463 => x"c178bff8",
   464 => x"c71ec01e",
   465 => x"87cafd49",
   466 => x"987086c8",
   467 => x"ff87ce02",
   468 => x"87c8fb49",
   469 => x"ff49dac1",
   470 => x"c187e9d7",
   471 => x"ebc5c34d",
   472 => x"c302bf97",
   473 => x"87ccd587",
   474 => x"bff0c5c3",
   475 => x"fbe5c24b",
   476 => x"ebc005bf",
   477 => x"49fdc387",
   478 => x"87c8d7ff",
   479 => x"ff49fac3",
   480 => x"7387c1d7",
   481 => x"99ffc349",
   482 => x"49c01e71",
   483 => x"7387c7fb",
   484 => x"29b7c849",
   485 => x"49c11e71",
   486 => x"c887fbfa",
   487 => x"87c1c686",
   488 => x"bff4c5c3",
   489 => x"dd029b4b",
   490 => x"f7e5c287",
   491 => x"dec749bf",
   492 => x"05987087",
   493 => x"4bc087c4",
   494 => x"e0c287d2",
   495 => x"87c3c749",
   496 => x"58fbe5c2",
   497 => x"e5c287c6",
   498 => x"78c048f7",
   499 => x"99c24973",
   500 => x"c387ce05",
   501 => x"d5ff49eb",
   502 => x"497087ea",
   503 => x"c20299c2",
   504 => x"734cfb87",
   505 => x"0599c149",
   506 => x"f4c387ce",
   507 => x"d3d5ff49",
   508 => x"c2497087",
   509 => x"87c20299",
   510 => x"49734cfa",
   511 => x"ce0599c8",
   512 => x"49f5c387",
   513 => x"87fcd4ff",
   514 => x"99c24970",
   515 => x"c387d502",
   516 => x"02bffcc5",
   517 => x"c14887ca",
   518 => x"c0c6c388",
   519 => x"87c2c058",
   520 => x"4dc14cff",
   521 => x"99c44973",
   522 => x"c387ce05",
   523 => x"d4ff49f2",
   524 => x"497087d2",
   525 => x"dc0299c2",
   526 => x"fcc5c387",
   527 => x"c7487ebf",
   528 => x"c003a8b7",
   529 => x"486e87cb",
   530 => x"c6c380c1",
   531 => x"c2c058c0",
   532 => x"c14cfe87",
   533 => x"49fdc34d",
   534 => x"87e8d3ff",
   535 => x"99c24970",
   536 => x"87d5c002",
   537 => x"bffcc5c3",
   538 => x"87c9c002",
   539 => x"48fcc5c3",
   540 => x"c2c078c0",
   541 => x"c14cfd87",
   542 => x"49fac34d",
   543 => x"87c4d3ff",
   544 => x"99c24970",
   545 => x"87d9c002",
   546 => x"bffcc5c3",
   547 => x"a8b7c748",
   548 => x"87c9c003",
   549 => x"48fcc5c3",
   550 => x"c2c078c7",
   551 => x"c14cfc87",
   552 => x"acb7c04d",
   553 => x"87d1c003",
   554 => x"c14a66c4",
   555 => x"026a82d8",
   556 => x"6a87c6c0",
   557 => x"7349744b",
   558 => x"c31ec00f",
   559 => x"dac11ef0",
   560 => x"87cef749",
   561 => x"987086c8",
   562 => x"87e2c002",
   563 => x"c348a6c8",
   564 => x"78bffcc5",
   565 => x"cb4966c8",
   566 => x"4866c491",
   567 => x"7e708071",
   568 => x"c002bf6e",
   569 => x"bf6e87c8",
   570 => x"4966c84b",
   571 => x"9d750f73",
   572 => x"87c8c002",
   573 => x"bffcc5c3",
   574 => x"87fbf249",
   575 => x"bfffe5c2",
   576 => x"87ddc002",
   577 => x"87c7c249",
   578 => x"c0029870",
   579 => x"c5c387d3",
   580 => x"f249bffc",
   581 => x"49c087e1",
   582 => x"c287c1f4",
   583 => x"c048ffe5",
   584 => x"f38ef478",
   585 => x"5e0e87db",
   586 => x"0e5d5c5b",
   587 => x"c34c711e",
   588 => x"49bff8c5",
   589 => x"4da1cdc1",
   590 => x"6981d1c1",
   591 => x"029c747e",
   592 => x"a5c487cf",
   593 => x"c37b744b",
   594 => x"49bff8c5",
   595 => x"6e87faf2",
   596 => x"059c747b",
   597 => x"4bc087c4",
   598 => x"4bc187c2",
   599 => x"fbf24973",
   600 => x"0266d487",
   601 => x"da4987c7",
   602 => x"c24a7087",
   603 => x"c24ac087",
   604 => x"265ac3e6",
   605 => x"0087caf2",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"1e000000",
   609 => x"c8ff4a71",
   610 => x"a17249bf",
   611 => x"1e4f2648",
   612 => x"89bfc8ff",
   613 => x"c0c0c0fe",
   614 => x"01a9c0c0",
   615 => x"4ac087c4",
   616 => x"4ac187c2",
   617 => x"4f264872",
   618 => x"5c5b5e0e",
   619 => x"4b710e5d",
   620 => x"d04cd4ff",
   621 => x"78c04866",
   622 => x"d8ff49d6",
   623 => x"ffc387cf",
   624 => x"c3496c7c",
   625 => x"4d7199ff",
   626 => x"99f0c349",
   627 => x"05a9e0c1",
   628 => x"ffc387cb",
   629 => x"c3486c7c",
   630 => x"0866d098",
   631 => x"7cffc378",
   632 => x"c8494a6c",
   633 => x"7cffc331",
   634 => x"b2714a6c",
   635 => x"31c84972",
   636 => x"6c7cffc3",
   637 => x"72b2714a",
   638 => x"c331c849",
   639 => x"4a6c7cff",
   640 => x"d0ffb271",
   641 => x"78e0c048",
   642 => x"c2029b73",
   643 => x"757b7287",
   644 => x"264d2648",
   645 => x"264b264c",
   646 => x"4f261e4f",
   647 => x"5c5b5e0e",
   648 => x"7686f80e",
   649 => x"49a6c81e",
   650 => x"c487fdfd",
   651 => x"6e4b7086",
   652 => x"03a8c248",
   653 => x"7387cac3",
   654 => x"9af0c34a",
   655 => x"02aad0c1",
   656 => x"e0c187c7",
   657 => x"f8c205aa",
   658 => x"c8497387",
   659 => x"87c30299",
   660 => x"7387c6ff",
   661 => x"c29cc34c",
   662 => x"cfc105ac",
   663 => x"4966c487",
   664 => x"1e7131c9",
   665 => x"c04a66c4",
   666 => x"c6c392f8",
   667 => x"817249c0",
   668 => x"87eac0fe",
   669 => x"1e4966c4",
   670 => x"ff49e3c0",
   671 => x"d887f3d5",
   672 => x"c8d5ff49",
   673 => x"1ec0c887",
   674 => x"49caf4c2",
   675 => x"87cbd9fd",
   676 => x"c048d0ff",
   677 => x"f4c278e0",
   678 => x"66d01eca",
   679 => x"92f8c04a",
   680 => x"49c0c6c3",
   681 => x"fbfd8172",
   682 => x"86d087f3",
   683 => x"c105acc1",
   684 => x"66c487cf",
   685 => x"7131c949",
   686 => x"4a66c41e",
   687 => x"c392f8c0",
   688 => x"7249c0c6",
   689 => x"d5fffd81",
   690 => x"caf4c287",
   691 => x"4a66c81e",
   692 => x"c392f8c0",
   693 => x"7249c0c6",
   694 => x"fdf9fd81",
   695 => x"4966c887",
   696 => x"49e3c01e",
   697 => x"87cad4ff",
   698 => x"d3ff49d7",
   699 => x"c0c887df",
   700 => x"caf4c21e",
   701 => x"ccd7fd49",
   702 => x"ff86d087",
   703 => x"e0c048d0",
   704 => x"fc8ef878",
   705 => x"5e0e87cd",
   706 => x"0e5d5c5b",
   707 => x"ff4d711e",
   708 => x"66d44cd4",
   709 => x"b7c3487e",
   710 => x"87c506a8",
   711 => x"e3c148c0",
   712 => x"fe497587",
   713 => x"7587efcf",
   714 => x"4b66c41e",
   715 => x"c393f8c0",
   716 => x"7383c0c6",
   717 => x"d4f4fd49",
   718 => x"6b83c887",
   719 => x"48d0ff4b",
   720 => x"dd78e1c8",
   721 => x"c349737c",
   722 => x"7c7199ff",
   723 => x"b7c84973",
   724 => x"99ffc329",
   725 => x"49737c71",
   726 => x"c329b7d0",
   727 => x"7c7199ff",
   728 => x"b7d84973",
   729 => x"c07c7129",
   730 => x"7c7c7c7c",
   731 => x"7c7c7c7c",
   732 => x"7c7c7c7c",
   733 => x"c478e0c0",
   734 => x"49dc1e66",
   735 => x"87f2d1ff",
   736 => x"487386c8",
   737 => x"87c9fa26",
   738 => x"5c5b5e0e",
   739 => x"711e0e5d",
   740 => x"4bd4ff7e",
   741 => x"c7c31e6e",
   742 => x"f2fd49f0",
   743 => x"86c487ef",
   744 => x"029d4d70",
   745 => x"c387c3c3",
   746 => x"4cbff8c7",
   747 => x"cdfe496e",
   748 => x"d0ff87e4",
   749 => x"78c5c848",
   750 => x"c07bd6c1",
   751 => x"c17b154a",
   752 => x"b7e0c082",
   753 => x"87f504aa",
   754 => x"c448d0ff",
   755 => x"78c5c878",
   756 => x"c17bd3c1",
   757 => x"7478c47b",
   758 => x"fcc1029c",
   759 => x"caf4c287",
   760 => x"4dc0c87e",
   761 => x"acb7c08c",
   762 => x"c887c603",
   763 => x"c04da4c0",
   764 => x"fbc0c34c",
   765 => x"d049bf97",
   766 => x"87d20299",
   767 => x"c7c31ec0",
   768 => x"f5fd49f0",
   769 => x"86c487d4",
   770 => x"c04a4970",
   771 => x"f4c287ef",
   772 => x"c7c31eca",
   773 => x"f5fd49f0",
   774 => x"86c487c0",
   775 => x"ff4a4970",
   776 => x"c5c848d0",
   777 => x"7bd4c178",
   778 => x"7bbf976e",
   779 => x"80c1486e",
   780 => x"8dc17e70",
   781 => x"87f0ff05",
   782 => x"c448d0ff",
   783 => x"059a7278",
   784 => x"48c087c5",
   785 => x"c187e5c0",
   786 => x"f0c7c31e",
   787 => x"e8f2fd49",
   788 => x"7486c487",
   789 => x"c4fe059c",
   790 => x"48d0ff87",
   791 => x"c178c5c8",
   792 => x"7bc07bd3",
   793 => x"48c178c4",
   794 => x"48c087c2",
   795 => x"264d2626",
   796 => x"264b264c",
   797 => x"5b5e0e4f",
   798 => x"4b710e5c",
   799 => x"d80266cc",
   800 => x"f0c04c87",
   801 => x"87d8028c",
   802 => x"8ac14a74",
   803 => x"8a87d102",
   804 => x"8a87cd02",
   805 => x"d787c902",
   806 => x"fb497387",
   807 => x"87d087ea",
   808 => x"49c01e74",
   809 => x"7487dff9",
   810 => x"f949731e",
   811 => x"86c887d8",
   812 => x"0087fcfe",
   813 => x"ddf3c21e",
   814 => x"b9c149bf",
   815 => x"59e1f3c2",
   816 => x"c348d4ff",
   817 => x"d0ff78ff",
   818 => x"78e1c848",
   819 => x"c148d4ff",
   820 => x"7131c478",
   821 => x"48d0ff78",
   822 => x"2678e0c0",
   823 => x"0000004f",
   824 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
