
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e8",x"c8",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"e8",x"c8",x"c3"),
    14 => (x"48",x"e4",x"f3",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c5",x"e2"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"e4",x"f3"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"f3",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"e4"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"e8",x"f3",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"ec",x"f3",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"ec",x"f3"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"f3",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"ec"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"f3",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"f3"),
   285 => (x"f3",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"f4"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"f5",x"f3",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"f5",x"f3",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"f6",x"f3"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"f3",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"f1"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"f2",x"f3"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"f3",x"f3",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"f4",x"f3"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"d2",x"fc",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"ca",x"f4"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"d0",x"f8",x"c0"),
   331 => (x"c0",x"f5",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f8",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"cc"),
   337 => (x"71",x"4a",x"dc",x"f5"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"d0",x"fb",x"c2",x"87"),
   343 => (x"fc",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"c8"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"d0",x"fb",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"ca",x"f4",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f8",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"cc"),
   359 => (x"71",x"4a",x"dc",x"f5"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"fc",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"d2"),
   364 => (x"f8",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"d0"),
   366 => (x"71",x"4a",x"c0",x"f5"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"c8",x"fc",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"c9",x"fc",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"ca",x"f4"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"d5",x"f4"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"f4",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"d6"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"d7",x"f4"),
   394 => (x"ce",x"fc",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"fc",x"c2",x"88",x"c1"),
   397 => (x"f4",x"c2",x"58",x"d2"),
   398 => (x"49",x"bf",x"97",x"d8"),
   399 => (x"f4",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"d9"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"df",x"c0",x"c3",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"da",x"f4"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"d2",x"fc",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"cc",x"f8",x"c0"),
   409 => (x"dc",x"f5",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"fc",x"c2",x"87",x"f8"),
   415 => (x"c3",x"4c",x"bf",x"ca"),
   416 => (x"c2",x"5c",x"f3",x"c0"),
   417 => (x"bf",x"97",x"ef",x"f4"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"ee",x"f4"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"f0",x"f4"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"f4",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"f1"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"df",x"c0",x"c3"),
   428 => (x"e7",x"c0",x"c3",x"81"),
   429 => (x"f7",x"f4",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"f6",x"f4",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"f8",x"f4",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"f9",x"f4",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"eb",x"c0",x"c3",x"4a"),
   440 => (x"e7",x"c0",x"c3",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"c0",x"c3",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"eb"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"dc",x"f4",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"db",x"f4",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"da",x"fc",x"c2"),
   450 => (x"bf",x"d6",x"fc",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"f3",x"c0",x"c3"),
   454 => (x"97",x"e1",x"f4",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"e0",x"f4",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"ef",x"c0",x"c3",x"82"),
   460 => (x"e7",x"c0",x"c3",x"5a"),
   461 => (x"c3",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"e3",x"c0"),
   463 => (x"c0",x"c3",x"78",x"a1"),
   464 => (x"c0",x"c3",x"48",x"f3"),
   465 => (x"c3",x"78",x"bf",x"e7"),
   466 => (x"c3",x"48",x"f7",x"c0"),
   467 => (x"78",x"bf",x"eb",x"c0"),
   468 => (x"bf",x"d2",x"fc",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"ef",x"c0",x"c3",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"fc",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"d6"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"d2",x"fc",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c3",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"df",x"c0"),
   489 => (x"bf",x"c8",x"f8",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"cc",x"f8",x"c0"),
   492 => (x"1e",x"ca",x"f4",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"d2",x"fc",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"ca",x"f4",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"f4",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"ca"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"d0",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"f2"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"da",x"fc"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"cf",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"f2"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"f8",x"0e",x"5d",x"5c"),
   533 => (x"9b",x"4b",x"71",x"86"),
   534 => (x"c0",x"87",x"c5",x"05"),
   535 => (x"87",x"d4",x"c2",x"48"),
   536 => (x"c0",x"4d",x"a3",x"c8"),
   537 => (x"02",x"66",x"d8",x"7d"),
   538 => (x"66",x"d8",x"87",x"c7"),
   539 => (x"c5",x"05",x"bf",x"97"),
   540 => (x"c1",x"48",x"c0",x"87"),
   541 => (x"66",x"d8",x"87",x"fe"),
   542 => (x"87",x"f2",x"fd",x"49"),
   543 => (x"02",x"6e",x"7e",x"70"),
   544 => (x"6e",x"87",x"ef",x"c1"),
   545 => (x"69",x"81",x"dc",x"49"),
   546 => (x"da",x"49",x"6e",x"7d"),
   547 => (x"4c",x"a3",x"c4",x"81"),
   548 => (x"c2",x"7c",x"69",x"9f"),
   549 => (x"02",x"bf",x"d2",x"fc"),
   550 => (x"49",x"6e",x"87",x"d0"),
   551 => (x"69",x"9f",x"81",x"d4"),
   552 => (x"ff",x"c0",x"4a",x"49"),
   553 => (x"32",x"d0",x"9a",x"ff"),
   554 => (x"4a",x"c0",x"87",x"c2"),
   555 => (x"6c",x"48",x"49",x"72"),
   556 => (x"c0",x"7c",x"70",x"80"),
   557 => (x"49",x"a3",x"cc",x"7b"),
   558 => (x"a3",x"d0",x"79",x"6c"),
   559 => (x"c4",x"79",x"c0",x"49"),
   560 => (x"78",x"c0",x"48",x"a6"),
   561 => (x"c4",x"4a",x"a3",x"d4"),
   562 => (x"91",x"c8",x"49",x"66"),
   563 => (x"c0",x"49",x"a1",x"72"),
   564 => (x"c4",x"79",x"6c",x"41"),
   565 => (x"80",x"c1",x"48",x"66"),
   566 => (x"c4",x"58",x"a6",x"c8"),
   567 => (x"ff",x"04",x"a8",x"b7"),
   568 => (x"4a",x"6d",x"87",x"e2"),
   569 => (x"2a",x"c5",x"2a",x"c9"),
   570 => (x"49",x"a3",x"f4",x"c0"),
   571 => (x"48",x"6e",x"79",x"72"),
   572 => (x"48",x"c0",x"87",x"c2"),
   573 => (x"fb",x"f9",x"8e",x"f8"),
   574 => (x"5b",x"5e",x"0e",x"87"),
   575 => (x"71",x"0e",x"5d",x"5c"),
   576 => (x"c8",x"f8",x"c0",x"4c"),
   577 => (x"74",x"78",x"ff",x"48"),
   578 => (x"ca",x"c1",x"02",x"9c"),
   579 => (x"49",x"a4",x"c8",x"87"),
   580 => (x"c2",x"c1",x"02",x"69"),
   581 => (x"4a",x"66",x"d0",x"87"),
   582 => (x"d4",x"82",x"49",x"6c"),
   583 => (x"66",x"d0",x"5a",x"a6"),
   584 => (x"fc",x"c2",x"b9",x"4d"),
   585 => (x"ff",x"4a",x"bf",x"ce"),
   586 => (x"71",x"99",x"72",x"ba"),
   587 => (x"e4",x"c0",x"02",x"99"),
   588 => (x"4b",x"a4",x"c4",x"87"),
   589 => (x"c3",x"f9",x"49",x"6b"),
   590 => (x"c2",x"7b",x"70",x"87"),
   591 => (x"49",x"bf",x"ca",x"fc"),
   592 => (x"7c",x"71",x"81",x"6c"),
   593 => (x"fc",x"c2",x"b9",x"75"),
   594 => (x"ff",x"4a",x"bf",x"ce"),
   595 => (x"71",x"99",x"72",x"ba"),
   596 => (x"dc",x"ff",x"05",x"99"),
   597 => (x"f8",x"7c",x"75",x"87"),
   598 => (x"73",x"1e",x"87",x"da"),
   599 => (x"9b",x"4b",x"71",x"1e"),
   600 => (x"c8",x"87",x"c7",x"02"),
   601 => (x"05",x"69",x"49",x"a3"),
   602 => (x"48",x"c0",x"87",x"c5"),
   603 => (x"c3",x"87",x"eb",x"c0"),
   604 => (x"4a",x"bf",x"e3",x"c0"),
   605 => (x"69",x"49",x"a3",x"c4"),
   606 => (x"c2",x"89",x"c2",x"49"),
   607 => (x"91",x"bf",x"ca",x"fc"),
   608 => (x"c2",x"4a",x"a2",x"71"),
   609 => (x"49",x"bf",x"ce",x"fc"),
   610 => (x"a2",x"71",x"99",x"6b"),
   611 => (x"1e",x"66",x"c8",x"4a"),
   612 => (x"e1",x"e9",x"49",x"72"),
   613 => (x"70",x"86",x"c4",x"87"),
   614 => (x"db",x"f7",x"48",x"49"),
   615 => (x"1e",x"73",x"1e",x"87"),
   616 => (x"02",x"9b",x"4b",x"71"),
   617 => (x"a3",x"c8",x"87",x"c7"),
   618 => (x"c5",x"05",x"69",x"49"),
   619 => (x"c0",x"48",x"c0",x"87"),
   620 => (x"c0",x"c3",x"87",x"eb"),
   621 => (x"c4",x"4a",x"bf",x"e3"),
   622 => (x"49",x"69",x"49",x"a3"),
   623 => (x"fc",x"c2",x"89",x"c2"),
   624 => (x"71",x"91",x"bf",x"ca"),
   625 => (x"fc",x"c2",x"4a",x"a2"),
   626 => (x"6b",x"49",x"bf",x"ce"),
   627 => (x"4a",x"a2",x"71",x"99"),
   628 => (x"72",x"1e",x"66",x"c8"),
   629 => (x"87",x"d4",x"e5",x"49"),
   630 => (x"49",x"70",x"86",x"c4"),
   631 => (x"87",x"d8",x"f6",x"48"),
   632 => (x"5c",x"5b",x"5e",x"0e"),
   633 => (x"86",x"f8",x"0e",x"5d"),
   634 => (x"a6",x"c4",x"4b",x"71"),
   635 => (x"c8",x"78",x"ff",x"48"),
   636 => (x"4d",x"69",x"49",x"a3"),
   637 => (x"a3",x"d4",x"4c",x"c0"),
   638 => (x"c8",x"49",x"74",x"4a"),
   639 => (x"49",x"a1",x"72",x"91"),
   640 => (x"66",x"d8",x"49",x"69"),
   641 => (x"70",x"88",x"71",x"48"),
   642 => (x"a9",x"66",x"d8",x"7e"),
   643 => (x"6e",x"87",x"ca",x"01"),
   644 => (x"87",x"c5",x"06",x"ad"),
   645 => (x"6e",x"5c",x"a6",x"c8"),
   646 => (x"c4",x"84",x"c1",x"4d"),
   647 => (x"ff",x"04",x"ac",x"b7"),
   648 => (x"48",x"66",x"87",x"d4"),
   649 => (x"cb",x"f5",x"8e",x"f8"),
   650 => (x"5b",x"5e",x"0e",x"87"),
   651 => (x"ec",x"0e",x"5d",x"5c"),
   652 => (x"59",x"a6",x"c8",x"86"),
   653 => (x"c1",x"48",x"a6",x"c8"),
   654 => (x"ff",x"ff",x"ff",x"ff"),
   655 => (x"80",x"c4",x"78",x"ff"),
   656 => (x"4d",x"c0",x"78",x"ff"),
   657 => (x"66",x"c4",x"4c",x"c0"),
   658 => (x"74",x"83",x"d4",x"4b"),
   659 => (x"73",x"91",x"c8",x"49"),
   660 => (x"4a",x"75",x"49",x"a1"),
   661 => (x"a2",x"73",x"92",x"c8"),
   662 => (x"6e",x"49",x"69",x"7e"),
   663 => (x"a6",x"d4",x"89",x"bf"),
   664 => (x"05",x"ad",x"74",x"59"),
   665 => (x"a6",x"d0",x"87",x"c6"),
   666 => (x"78",x"bf",x"6e",x"48"),
   667 => (x"c0",x"48",x"66",x"d0"),
   668 => (x"cf",x"04",x"a8",x"b7"),
   669 => (x"49",x"66",x"d0",x"87"),
   670 => (x"03",x"a9",x"66",x"c8"),
   671 => (x"a6",x"d0",x"87",x"c6"),
   672 => (x"59",x"a6",x"cc",x"5c"),
   673 => (x"b7",x"c4",x"84",x"c1"),
   674 => (x"f9",x"fe",x"04",x"ac"),
   675 => (x"c4",x"85",x"c1",x"87"),
   676 => (x"fe",x"04",x"ad",x"b7"),
   677 => (x"66",x"cc",x"87",x"ee"),
   678 => (x"f3",x"8e",x"ec",x"48"),
   679 => (x"5e",x"0e",x"87",x"d6"),
   680 => (x"0e",x"5d",x"5c",x"5b"),
   681 => (x"4b",x"71",x"86",x"f0"),
   682 => (x"4c",x"66",x"e0",x"c0"),
   683 => (x"9b",x"73",x"2c",x"c9"),
   684 => (x"87",x"e1",x"c3",x"02"),
   685 => (x"69",x"49",x"a3",x"c8"),
   686 => (x"87",x"d9",x"c3",x"02"),
   687 => (x"c0",x"49",x"a3",x"d0"),
   688 => (x"6b",x"79",x"66",x"e0"),
   689 => (x"c3",x"02",x"ac",x"7e"),
   690 => (x"fc",x"c2",x"87",x"cb"),
   691 => (x"ff",x"49",x"bf",x"ce"),
   692 => (x"74",x"4a",x"71",x"b9"),
   693 => (x"6e",x"48",x"71",x"9a"),
   694 => (x"58",x"a6",x"cc",x"98"),
   695 => (x"c4",x"4d",x"a3",x"c4"),
   696 => (x"78",x"6d",x"48",x"a6"),
   697 => (x"05",x"aa",x"66",x"c8"),
   698 => (x"7b",x"74",x"87",x"c5"),
   699 => (x"72",x"87",x"d1",x"c2"),
   700 => (x"fb",x"49",x"73",x"1e"),
   701 => (x"86",x"c4",x"87",x"ea"),
   702 => (x"c0",x"48",x"7e",x"70"),
   703 => (x"d0",x"04",x"a8",x"b7"),
   704 => (x"4a",x"a3",x"d4",x"87"),
   705 => (x"91",x"c8",x"49",x"6e"),
   706 => (x"21",x"49",x"a1",x"72"),
   707 => (x"c7",x"7d",x"69",x"7b"),
   708 => (x"cc",x"7b",x"c0",x"87"),
   709 => (x"7d",x"69",x"49",x"a3"),
   710 => (x"73",x"1e",x"66",x"c8"),
   711 => (x"87",x"c0",x"fb",x"49"),
   712 => (x"7e",x"70",x"86",x"c4"),
   713 => (x"49",x"a3",x"f4",x"c0"),
   714 => (x"69",x"48",x"a6",x"cc"),
   715 => (x"48",x"66",x"c8",x"78"),
   716 => (x"06",x"a8",x"66",x"cc"),
   717 => (x"48",x"6e",x"87",x"c9"),
   718 => (x"04",x"a8",x"b7",x"c0"),
   719 => (x"6e",x"87",x"e0",x"c0"),
   720 => (x"a8",x"b7",x"c0",x"48"),
   721 => (x"87",x"ec",x"c0",x"04"),
   722 => (x"6e",x"4a",x"a3",x"d4"),
   723 => (x"72",x"91",x"c8",x"49"),
   724 => (x"66",x"c8",x"49",x"a1"),
   725 => (x"70",x"88",x"69",x"48"),
   726 => (x"a9",x"66",x"cc",x"49"),
   727 => (x"73",x"87",x"d5",x"06"),
   728 => (x"87",x"c5",x"fb",x"49"),
   729 => (x"a3",x"d4",x"49",x"70"),
   730 => (x"72",x"91",x"c8",x"4a"),
   731 => (x"66",x"c8",x"49",x"a1"),
   732 => (x"79",x"66",x"c4",x"41"),
   733 => (x"49",x"74",x"8c",x"6b"),
   734 => (x"f5",x"49",x"73",x"1e"),
   735 => (x"86",x"c4",x"87",x"fb"),
   736 => (x"49",x"66",x"e0",x"c0"),
   737 => (x"02",x"99",x"ff",x"c7"),
   738 => (x"f4",x"c2",x"87",x"cb"),
   739 => (x"49",x"73",x"1e",x"ca"),
   740 => (x"c4",x"87",x"c7",x"f7"),
   741 => (x"ef",x"8e",x"f0",x"86"),
   742 => (x"73",x"1e",x"87",x"da"),
   743 => (x"9b",x"4b",x"71",x"1e"),
   744 => (x"87",x"e4",x"c0",x"02"),
   745 => (x"5b",x"f7",x"c0",x"c3"),
   746 => (x"8a",x"c2",x"4a",x"73"),
   747 => (x"bf",x"ca",x"fc",x"c2"),
   748 => (x"c0",x"c3",x"92",x"49"),
   749 => (x"72",x"48",x"bf",x"e3"),
   750 => (x"fb",x"c0",x"c3",x"80"),
   751 => (x"c4",x"48",x"71",x"58"),
   752 => (x"da",x"fc",x"c2",x"30"),
   753 => (x"87",x"ed",x"c0",x"58"),
   754 => (x"48",x"f3",x"c0",x"c3"),
   755 => (x"bf",x"e7",x"c0",x"c3"),
   756 => (x"f7",x"c0",x"c3",x"78"),
   757 => (x"eb",x"c0",x"c3",x"48"),
   758 => (x"fc",x"c2",x"78",x"bf"),
   759 => (x"c9",x"02",x"bf",x"d2"),
   760 => (x"ca",x"fc",x"c2",x"87"),
   761 => (x"31",x"c4",x"49",x"bf"),
   762 => (x"c0",x"c3",x"87",x"c7"),
   763 => (x"c4",x"49",x"bf",x"ef"),
   764 => (x"da",x"fc",x"c2",x"31"),
   765 => (x"87",x"c0",x"ee",x"59"),
   766 => (x"5c",x"5b",x"5e",x"0e"),
   767 => (x"c0",x"4a",x"71",x"0e"),
   768 => (x"02",x"9a",x"72",x"4b"),
   769 => (x"da",x"87",x"e1",x"c0"),
   770 => (x"69",x"9f",x"49",x"a2"),
   771 => (x"d2",x"fc",x"c2",x"4b"),
   772 => (x"87",x"cf",x"02",x"bf"),
   773 => (x"9f",x"49",x"a2",x"d4"),
   774 => (x"c0",x"4c",x"49",x"69"),
   775 => (x"d0",x"9c",x"ff",x"ff"),
   776 => (x"c0",x"87",x"c2",x"34"),
   777 => (x"b3",x"49",x"74",x"4c"),
   778 => (x"ed",x"fd",x"49",x"73"),
   779 => (x"87",x"c6",x"ed",x"87"),
   780 => (x"5c",x"5b",x"5e",x"0e"),
   781 => (x"86",x"f4",x"0e",x"5d"),
   782 => (x"7e",x"c0",x"4a",x"71"),
   783 => (x"d8",x"02",x"9a",x"72"),
   784 => (x"c6",x"f4",x"c2",x"87"),
   785 => (x"c2",x"78",x"c0",x"48"),
   786 => (x"c3",x"48",x"fe",x"f3"),
   787 => (x"78",x"bf",x"f7",x"c0"),
   788 => (x"48",x"c2",x"f4",x"c2"),
   789 => (x"bf",x"f3",x"c0",x"c3"),
   790 => (x"e7",x"fc",x"c2",x"78"),
   791 => (x"c2",x"50",x"c0",x"48"),
   792 => (x"49",x"bf",x"d6",x"fc"),
   793 => (x"bf",x"c6",x"f4",x"c2"),
   794 => (x"03",x"aa",x"71",x"4a"),
   795 => (x"72",x"87",x"c0",x"c4"),
   796 => (x"05",x"99",x"cf",x"49"),
   797 => (x"c2",x"87",x"e1",x"c0"),
   798 => (x"c2",x"1e",x"ca",x"f4"),
   799 => (x"49",x"bf",x"fe",x"f3"),
   800 => (x"48",x"fe",x"f3",x"c2"),
   801 => (x"71",x"78",x"a1",x"c1"),
   802 => (x"87",x"ea",x"dd",x"ff"),
   803 => (x"f8",x"c0",x"86",x"c4"),
   804 => (x"f4",x"c2",x"48",x"c4"),
   805 => (x"87",x"cc",x"78",x"ca"),
   806 => (x"bf",x"c4",x"f8",x"c0"),
   807 => (x"80",x"e0",x"c0",x"48"),
   808 => (x"58",x"c8",x"f8",x"c0"),
   809 => (x"bf",x"c6",x"f4",x"c2"),
   810 => (x"c2",x"80",x"c1",x"48"),
   811 => (x"27",x"58",x"ca",x"f4"),
   812 => (x"00",x"00",x"0e",x"04"),
   813 => (x"4d",x"bf",x"97",x"bf"),
   814 => (x"e2",x"c2",x"02",x"9d"),
   815 => (x"ad",x"e5",x"c3",x"87"),
   816 => (x"87",x"db",x"c2",x"02"),
   817 => (x"bf",x"c4",x"f8",x"c0"),
   818 => (x"49",x"a3",x"cb",x"4b"),
   819 => (x"ac",x"cf",x"4c",x"11"),
   820 => (x"87",x"d2",x"c1",x"05"),
   821 => (x"99",x"df",x"49",x"75"),
   822 => (x"91",x"cd",x"89",x"c1"),
   823 => (x"81",x"da",x"fc",x"c2"),
   824 => (x"12",x"4a",x"a3",x"c1"),
   825 => (x"4a",x"a3",x"c3",x"51"),
   826 => (x"a3",x"c5",x"51",x"12"),
   827 => (x"c7",x"51",x"12",x"4a"),
   828 => (x"51",x"12",x"4a",x"a3"),
   829 => (x"12",x"4a",x"a3",x"c9"),
   830 => (x"4a",x"a3",x"ce",x"51"),
   831 => (x"a3",x"d0",x"51",x"12"),
   832 => (x"d2",x"51",x"12",x"4a"),
   833 => (x"51",x"12",x"4a",x"a3"),
   834 => (x"12",x"4a",x"a3",x"d4"),
   835 => (x"4a",x"a3",x"d6",x"51"),
   836 => (x"a3",x"d8",x"51",x"12"),
   837 => (x"dc",x"51",x"12",x"4a"),
   838 => (x"51",x"12",x"4a",x"a3"),
   839 => (x"12",x"4a",x"a3",x"de"),
   840 => (x"c0",x"7e",x"c1",x"51"),
   841 => (x"49",x"74",x"87",x"f9"),
   842 => (x"c0",x"05",x"99",x"c8"),
   843 => (x"49",x"74",x"87",x"ea"),
   844 => (x"d0",x"05",x"99",x"d0"),
   845 => (x"02",x"66",x"dc",x"87"),
   846 => (x"73",x"87",x"ca",x"c0"),
   847 => (x"0f",x"66",x"dc",x"49"),
   848 => (x"d3",x"02",x"98",x"70"),
   849 => (x"c0",x"05",x"6e",x"87"),
   850 => (x"fc",x"c2",x"87",x"c6"),
   851 => (x"50",x"c0",x"48",x"da"),
   852 => (x"bf",x"c4",x"f8",x"c0"),
   853 => (x"87",x"e7",x"c2",x"48"),
   854 => (x"48",x"e7",x"fc",x"c2"),
   855 => (x"c2",x"7e",x"50",x"c0"),
   856 => (x"49",x"bf",x"d6",x"fc"),
   857 => (x"bf",x"c6",x"f4",x"c2"),
   858 => (x"04",x"aa",x"71",x"4a"),
   859 => (x"c3",x"87",x"c0",x"fc"),
   860 => (x"05",x"bf",x"f7",x"c0"),
   861 => (x"c2",x"87",x"c8",x"c0"),
   862 => (x"02",x"bf",x"d2",x"fc"),
   863 => (x"c0",x"87",x"fe",x"c1"),
   864 => (x"ff",x"48",x"c8",x"f8"),
   865 => (x"c2",x"f4",x"c2",x"78"),
   866 => (x"ef",x"e7",x"49",x"bf"),
   867 => (x"c2",x"49",x"70",x"87"),
   868 => (x"c4",x"59",x"c6",x"f4"),
   869 => (x"f4",x"c2",x"48",x"a6"),
   870 => (x"c2",x"78",x"bf",x"c2"),
   871 => (x"02",x"bf",x"d2",x"fc"),
   872 => (x"c4",x"87",x"d8",x"c0"),
   873 => (x"ff",x"cf",x"49",x"66"),
   874 => (x"99",x"f8",x"ff",x"ff"),
   875 => (x"c5",x"c0",x"02",x"a9"),
   876 => (x"c0",x"4d",x"c0",x"87"),
   877 => (x"4d",x"c1",x"87",x"e1"),
   878 => (x"c4",x"87",x"dc",x"c0"),
   879 => (x"ff",x"cf",x"49",x"66"),
   880 => (x"02",x"a9",x"99",x"f8"),
   881 => (x"c8",x"87",x"c8",x"c0"),
   882 => (x"78",x"c0",x"48",x"a6"),
   883 => (x"c8",x"87",x"c5",x"c0"),
   884 => (x"78",x"c1",x"48",x"a6"),
   885 => (x"75",x"4d",x"66",x"c8"),
   886 => (x"e0",x"c0",x"05",x"9d"),
   887 => (x"49",x"66",x"c4",x"87"),
   888 => (x"fc",x"c2",x"89",x"c2"),
   889 => (x"91",x"4a",x"bf",x"ca"),
   890 => (x"bf",x"e3",x"c0",x"c3"),
   891 => (x"fe",x"f3",x"c2",x"4a"),
   892 => (x"78",x"a1",x"72",x"48"),
   893 => (x"48",x"c6",x"f4",x"c2"),
   894 => (x"e2",x"f9",x"78",x"c0"),
   895 => (x"f4",x"48",x"c0",x"87"),
   896 => (x"87",x"f0",x"e5",x"8e"),
   897 => (x"00",x"00",x"00",x"00"),
   898 => (x"ff",x"ff",x"ff",x"ff"),
   899 => (x"00",x"00",x"0e",x"14"),
   900 => (x"00",x"00",x"0e",x"1d"),
   901 => (x"33",x"54",x"41",x"46"),
   902 => (x"20",x"20",x"20",x"32"),
   903 => (x"54",x"41",x"46",x"00"),
   904 => (x"20",x"20",x"36",x"31"),
   905 => (x"ff",x"1e",x"00",x"20"),
   906 => (x"ff",x"c3",x"48",x"d4"),
   907 => (x"26",x"48",x"68",x"78"),
   908 => (x"d4",x"ff",x"1e",x"4f"),
   909 => (x"78",x"ff",x"c3",x"48"),
   910 => (x"c8",x"48",x"d0",x"ff"),
   911 => (x"d4",x"ff",x"78",x"e1"),
   912 => (x"c3",x"78",x"d4",x"48"),
   913 => (x"ff",x"48",x"fb",x"c0"),
   914 => (x"26",x"50",x"bf",x"d4"),
   915 => (x"d0",x"ff",x"1e",x"4f"),
   916 => (x"78",x"e0",x"c0",x"48"),
   917 => (x"ff",x"1e",x"4f",x"26"),
   918 => (x"49",x"70",x"87",x"cc"),
   919 => (x"87",x"c6",x"02",x"99"),
   920 => (x"05",x"a9",x"fb",x"c0"),
   921 => (x"48",x"71",x"87",x"f1"),
   922 => (x"5e",x"0e",x"4f",x"26"),
   923 => (x"71",x"0e",x"5c",x"5b"),
   924 => (x"fe",x"4c",x"c0",x"4b"),
   925 => (x"49",x"70",x"87",x"f0"),
   926 => (x"f9",x"c0",x"02",x"99"),
   927 => (x"a9",x"ec",x"c0",x"87"),
   928 => (x"87",x"f2",x"c0",x"02"),
   929 => (x"02",x"a9",x"fb",x"c0"),
   930 => (x"cc",x"87",x"eb",x"c0"),
   931 => (x"03",x"ac",x"b7",x"66"),
   932 => (x"66",x"d0",x"87",x"c7"),
   933 => (x"71",x"87",x"c2",x"02"),
   934 => (x"02",x"99",x"71",x"53"),
   935 => (x"84",x"c1",x"87",x"c2"),
   936 => (x"70",x"87",x"c3",x"fe"),
   937 => (x"cd",x"02",x"99",x"49"),
   938 => (x"a9",x"ec",x"c0",x"87"),
   939 => (x"c0",x"87",x"c7",x"02"),
   940 => (x"ff",x"05",x"a9",x"fb"),
   941 => (x"66",x"d0",x"87",x"d5"),
   942 => (x"c0",x"87",x"c3",x"02"),
   943 => (x"ec",x"c0",x"7b",x"97"),
   944 => (x"87",x"c4",x"05",x"a9"),
   945 => (x"87",x"c5",x"4a",x"74"),
   946 => (x"0a",x"c0",x"4a",x"74"),
   947 => (x"c2",x"48",x"72",x"8a"),
   948 => (x"26",x"4d",x"26",x"87"),
   949 => (x"26",x"4b",x"26",x"4c"),
   950 => (x"c9",x"fd",x"1e",x"4f"),
   951 => (x"c0",x"49",x"70",x"87"),
   952 => (x"04",x"a9",x"b7",x"f0"),
   953 => (x"f9",x"c0",x"87",x"ca"),
   954 => (x"c3",x"01",x"a9",x"b7"),
   955 => (x"89",x"f0",x"c0",x"87"),
   956 => (x"a9",x"b7",x"c1",x"c1"),
   957 => (x"c1",x"87",x"ca",x"04"),
   958 => (x"01",x"a9",x"b7",x"da"),
   959 => (x"f7",x"c0",x"87",x"c3"),
   960 => (x"b7",x"e1",x"c1",x"89"),
   961 => (x"87",x"ca",x"04",x"a9"),
   962 => (x"a9",x"b7",x"fa",x"c1"),
   963 => (x"c0",x"87",x"c3",x"01"),
   964 => (x"48",x"71",x"89",x"fd"),
   965 => (x"5e",x"0e",x"4f",x"26"),
   966 => (x"71",x"0e",x"5c",x"5b"),
   967 => (x"4c",x"d4",x"ff",x"4a"),
   968 => (x"ea",x"c0",x"49",x"72"),
   969 => (x"9b",x"4b",x"70",x"87"),
   970 => (x"c1",x"87",x"c2",x"02"),
   971 => (x"48",x"d0",x"ff",x"8b"),
   972 => (x"c1",x"78",x"c5",x"c8"),
   973 => (x"49",x"73",x"7c",x"d5"),
   974 => (x"f2",x"c2",x"31",x"c6"),
   975 => (x"4a",x"bf",x"97",x"f3"),
   976 => (x"70",x"b0",x"71",x"48"),
   977 => (x"48",x"d0",x"ff",x"7c"),
   978 => (x"48",x"73",x"78",x"c4"),
   979 => (x"0e",x"87",x"c4",x"fe"),
   980 => (x"5d",x"5c",x"5b",x"5e"),
   981 => (x"71",x"86",x"f8",x"0e"),
   982 => (x"fb",x"7e",x"c0",x"4c"),
   983 => (x"4b",x"c0",x"87",x"d3"),
   984 => (x"97",x"fc",x"ff",x"c0"),
   985 => (x"a9",x"c0",x"49",x"bf"),
   986 => (x"fb",x"87",x"cf",x"04"),
   987 => (x"83",x"c1",x"87",x"e8"),
   988 => (x"97",x"fc",x"ff",x"c0"),
   989 => (x"06",x"ab",x"49",x"bf"),
   990 => (x"ff",x"c0",x"87",x"f1"),
   991 => (x"02",x"bf",x"97",x"fc"),
   992 => (x"e1",x"fa",x"87",x"cf"),
   993 => (x"99",x"49",x"70",x"87"),
   994 => (x"c0",x"87",x"c6",x"02"),
   995 => (x"f1",x"05",x"a9",x"ec"),
   996 => (x"fa",x"4b",x"c0",x"87"),
   997 => (x"4d",x"70",x"87",x"d0"),
   998 => (x"c8",x"87",x"cb",x"fa"),
   999 => (x"c5",x"fa",x"58",x"a6"),
  1000 => (x"c1",x"4a",x"70",x"87"),
  1001 => (x"49",x"a4",x"c8",x"83"),
  1002 => (x"ad",x"49",x"69",x"97"),
  1003 => (x"c0",x"87",x"c7",x"02"),
  1004 => (x"c0",x"05",x"ad",x"ff"),
  1005 => (x"a4",x"c9",x"87",x"e7"),
  1006 => (x"49",x"69",x"97",x"49"),
  1007 => (x"02",x"a9",x"66",x"c4"),
  1008 => (x"c0",x"48",x"87",x"c7"),
  1009 => (x"d4",x"05",x"a8",x"ff"),
  1010 => (x"49",x"a4",x"ca",x"87"),
  1011 => (x"aa",x"49",x"69",x"97"),
  1012 => (x"c0",x"87",x"c6",x"02"),
  1013 => (x"c4",x"05",x"aa",x"ff"),
  1014 => (x"d0",x"7e",x"c1",x"87"),
  1015 => (x"ad",x"ec",x"c0",x"87"),
  1016 => (x"c0",x"87",x"c6",x"02"),
  1017 => (x"c4",x"05",x"ad",x"fb"),
  1018 => (x"c1",x"4b",x"c0",x"87"),
  1019 => (x"fe",x"02",x"6e",x"7e"),
  1020 => (x"d8",x"f9",x"87",x"e1"),
  1021 => (x"f8",x"48",x"73",x"87"),
  1022 => (x"87",x"d5",x"fb",x"8e"),
  1023 => (x"5b",x"5e",x"0e",x"00"),
  1024 => (x"1e",x"0e",x"5d",x"5c"),
  1025 => (x"4c",x"c0",x"4b",x"71"),
  1026 => (x"c0",x"04",x"ab",x"4d"),
  1027 => (x"fd",x"c0",x"87",x"e8"),
  1028 => (x"9d",x"75",x"1e",x"cf"),
  1029 => (x"c0",x"87",x"c4",x"02"),
  1030 => (x"c1",x"87",x"c2",x"4a"),
  1031 => (x"f0",x"49",x"72",x"4a"),
  1032 => (x"86",x"c4",x"87",x"ce"),
  1033 => (x"84",x"c1",x"7e",x"70"),
  1034 => (x"87",x"c2",x"05",x"6e"),
  1035 => (x"85",x"c1",x"4c",x"73"),
  1036 => (x"ff",x"06",x"ac",x"73"),
  1037 => (x"48",x"6e",x"87",x"d8"),
  1038 => (x"26",x"4d",x"26",x"26"),
  1039 => (x"26",x"4b",x"26",x"4c"),
  1040 => (x"5b",x"5e",x"0e",x"4f"),
  1041 => (x"1e",x"0e",x"5d",x"5c"),
  1042 => (x"de",x"49",x"4c",x"71"),
  1043 => (x"d5",x"c1",x"c3",x"91"),
  1044 => (x"97",x"85",x"71",x"4d"),
  1045 => (x"dd",x"c1",x"02",x"6d"),
  1046 => (x"c0",x"c1",x"c3",x"87"),
  1047 => (x"82",x"74",x"4a",x"bf"),
  1048 => (x"d8",x"fe",x"49",x"72"),
  1049 => (x"6e",x"7e",x"70",x"87"),
  1050 => (x"87",x"f3",x"c0",x"02"),
  1051 => (x"4b",x"c8",x"c1",x"c3"),
  1052 => (x"49",x"cb",x"4a",x"6e"),
  1053 => (x"87",x"f0",x"c0",x"ff"),
  1054 => (x"93",x"cb",x"4b",x"74"),
  1055 => (x"83",x"f5",x"e3",x"c1"),
  1056 => (x"c2",x"c1",x"83",x"c4"),
  1057 => (x"49",x"74",x"7b",x"fa"),
  1058 => (x"87",x"eb",x"d4",x"c1"),
  1059 => (x"c1",x"c3",x"7b",x"75"),
  1060 => (x"49",x"bf",x"97",x"d4"),
  1061 => (x"c8",x"c1",x"c3",x"1e"),
  1062 => (x"d8",x"ef",x"c1",x"49"),
  1063 => (x"74",x"86",x"c4",x"87"),
  1064 => (x"d2",x"d4",x"c1",x"49"),
  1065 => (x"c1",x"49",x"c0",x"87"),
  1066 => (x"c3",x"87",x"f1",x"d5"),
  1067 => (x"c0",x"48",x"fc",x"c0"),
  1068 => (x"dd",x"49",x"c1",x"78"),
  1069 => (x"fd",x"26",x"87",x"d0"),
  1070 => (x"6f",x"4c",x"87",x"ff"),
  1071 => (x"6e",x"69",x"64",x"61"),
  1072 => (x"2e",x"2e",x"2e",x"67"),
  1073 => (x"5b",x"5e",x"0e",x"00"),
  1074 => (x"4b",x"71",x"0e",x"5c"),
  1075 => (x"c0",x"c1",x"c3",x"4a"),
  1076 => (x"49",x"72",x"82",x"bf"),
  1077 => (x"70",x"87",x"e6",x"fc"),
  1078 => (x"c4",x"02",x"9c",x"4c"),
  1079 => (x"d7",x"ec",x"49",x"87"),
  1080 => (x"c0",x"c1",x"c3",x"87"),
  1081 => (x"c1",x"78",x"c0",x"48"),
  1082 => (x"87",x"da",x"dc",x"49"),
  1083 => (x"0e",x"87",x"cc",x"fd"),
  1084 => (x"5d",x"5c",x"5b",x"5e"),
  1085 => (x"c2",x"86",x"f4",x"0e"),
  1086 => (x"c0",x"4d",x"ca",x"f4"),
  1087 => (x"48",x"a6",x"c4",x"4c"),
  1088 => (x"c1",x"c3",x"78",x"c0"),
  1089 => (x"c0",x"49",x"bf",x"c0"),
  1090 => (x"c1",x"c1",x"06",x"a9"),
  1091 => (x"ca",x"f4",x"c2",x"87"),
  1092 => (x"c0",x"02",x"98",x"48"),
  1093 => (x"fd",x"c0",x"87",x"f8"),
  1094 => (x"66",x"c8",x"1e",x"cf"),
  1095 => (x"c4",x"87",x"c7",x"02"),
  1096 => (x"78",x"c0",x"48",x"a6"),
  1097 => (x"a6",x"c4",x"87",x"c5"),
  1098 => (x"c4",x"78",x"c1",x"48"),
  1099 => (x"ff",x"eb",x"49",x"66"),
  1100 => (x"70",x"86",x"c4",x"87"),
  1101 => (x"c4",x"84",x"c1",x"4d"),
  1102 => (x"80",x"c1",x"48",x"66"),
  1103 => (x"c3",x"58",x"a6",x"c8"),
  1104 => (x"49",x"bf",x"c0",x"c1"),
  1105 => (x"87",x"c6",x"03",x"ac"),
  1106 => (x"ff",x"05",x"9d",x"75"),
  1107 => (x"4c",x"c0",x"87",x"c8"),
  1108 => (x"c3",x"02",x"9d",x"75"),
  1109 => (x"fd",x"c0",x"87",x"e0"),
  1110 => (x"66",x"c8",x"1e",x"cf"),
  1111 => (x"cc",x"87",x"c7",x"02"),
  1112 => (x"78",x"c0",x"48",x"a6"),
  1113 => (x"a6",x"cc",x"87",x"c5"),
  1114 => (x"cc",x"78",x"c1",x"48"),
  1115 => (x"ff",x"ea",x"49",x"66"),
  1116 => (x"70",x"86",x"c4",x"87"),
  1117 => (x"c2",x"02",x"6e",x"7e"),
  1118 => (x"49",x"6e",x"87",x"e9"),
  1119 => (x"69",x"97",x"81",x"cb"),
  1120 => (x"02",x"99",x"d0",x"49"),
  1121 => (x"c1",x"87",x"d6",x"c1"),
  1122 => (x"74",x"4a",x"c5",x"c3"),
  1123 => (x"c1",x"91",x"cb",x"49"),
  1124 => (x"72",x"81",x"f5",x"e3"),
  1125 => (x"c3",x"81",x"c8",x"79"),
  1126 => (x"49",x"74",x"51",x"ff"),
  1127 => (x"c1",x"c3",x"91",x"de"),
  1128 => (x"85",x"71",x"4d",x"d5"),
  1129 => (x"7d",x"97",x"c1",x"c2"),
  1130 => (x"c0",x"49",x"a5",x"c1"),
  1131 => (x"fc",x"c2",x"51",x"e0"),
  1132 => (x"02",x"bf",x"97",x"da"),
  1133 => (x"84",x"c1",x"87",x"d2"),
  1134 => (x"c2",x"4b",x"a5",x"c2"),
  1135 => (x"db",x"4a",x"da",x"fc"),
  1136 => (x"e3",x"fb",x"fe",x"49"),
  1137 => (x"87",x"db",x"c1",x"87"),
  1138 => (x"c0",x"49",x"a5",x"cd"),
  1139 => (x"c2",x"84",x"c1",x"51"),
  1140 => (x"4a",x"6e",x"4b",x"a5"),
  1141 => (x"fb",x"fe",x"49",x"cb"),
  1142 => (x"c6",x"c1",x"87",x"ce"),
  1143 => (x"c1",x"c1",x"c1",x"87"),
  1144 => (x"cb",x"49",x"74",x"4a"),
  1145 => (x"f5",x"e3",x"c1",x"91"),
  1146 => (x"c2",x"79",x"72",x"81"),
  1147 => (x"bf",x"97",x"da",x"fc"),
  1148 => (x"74",x"87",x"d8",x"02"),
  1149 => (x"c1",x"91",x"de",x"49"),
  1150 => (x"d5",x"c1",x"c3",x"84"),
  1151 => (x"c2",x"83",x"71",x"4b"),
  1152 => (x"dd",x"4a",x"da",x"fc"),
  1153 => (x"df",x"fa",x"fe",x"49"),
  1154 => (x"74",x"87",x"d8",x"87"),
  1155 => (x"c3",x"93",x"de",x"4b"),
  1156 => (x"cb",x"83",x"d5",x"c1"),
  1157 => (x"51",x"c0",x"49",x"a3"),
  1158 => (x"6e",x"73",x"84",x"c1"),
  1159 => (x"fe",x"49",x"cb",x"4a"),
  1160 => (x"c4",x"87",x"c5",x"fa"),
  1161 => (x"80",x"c1",x"48",x"66"),
  1162 => (x"c7",x"58",x"a6",x"c8"),
  1163 => (x"c5",x"c0",x"03",x"ac"),
  1164 => (x"fc",x"05",x"6e",x"87"),
  1165 => (x"48",x"74",x"87",x"e0"),
  1166 => (x"fc",x"f7",x"8e",x"f4"),
  1167 => (x"1e",x"73",x"1e",x"87"),
  1168 => (x"cb",x"49",x"4b",x"71"),
  1169 => (x"f5",x"e3",x"c1",x"91"),
  1170 => (x"4a",x"a1",x"c8",x"81"),
  1171 => (x"48",x"f3",x"f2",x"c2"),
  1172 => (x"a1",x"c9",x"50",x"12"),
  1173 => (x"fc",x"ff",x"c0",x"4a"),
  1174 => (x"ca",x"50",x"12",x"48"),
  1175 => (x"d4",x"c1",x"c3",x"81"),
  1176 => (x"c3",x"50",x"11",x"48"),
  1177 => (x"bf",x"97",x"d4",x"c1"),
  1178 => (x"49",x"c0",x"1e",x"49"),
  1179 => (x"87",x"c5",x"e8",x"c1"),
  1180 => (x"48",x"fc",x"c0",x"c3"),
  1181 => (x"49",x"c1",x"78",x"de"),
  1182 => (x"26",x"87",x"cb",x"d6"),
  1183 => (x"1e",x"87",x"fe",x"f6"),
  1184 => (x"cb",x"49",x"4a",x"71"),
  1185 => (x"f5",x"e3",x"c1",x"91"),
  1186 => (x"11",x"81",x"c8",x"81"),
  1187 => (x"c0",x"c1",x"c3",x"48"),
  1188 => (x"c0",x"c1",x"c3",x"58"),
  1189 => (x"c1",x"78",x"c0",x"48"),
  1190 => (x"87",x"ea",x"d5",x"49"),
  1191 => (x"c0",x"1e",x"4f",x"26"),
  1192 => (x"f7",x"cd",x"c1",x"49"),
  1193 => (x"1e",x"4f",x"26",x"87"),
  1194 => (x"d2",x"02",x"99",x"71"),
  1195 => (x"ca",x"e5",x"c1",x"87"),
  1196 => (x"f7",x"50",x"c0",x"48"),
  1197 => (x"ff",x"c9",x"c1",x"80"),
  1198 => (x"ee",x"e3",x"c1",x"40"),
  1199 => (x"c1",x"87",x"ce",x"78"),
  1200 => (x"c1",x"48",x"c6",x"e5"),
  1201 => (x"fc",x"78",x"e7",x"e3"),
  1202 => (x"de",x"ca",x"c1",x"80"),
  1203 => (x"0e",x"4f",x"26",x"78"),
  1204 => (x"0e",x"5c",x"5b",x"5e"),
  1205 => (x"cb",x"4a",x"4c",x"71"),
  1206 => (x"f5",x"e3",x"c1",x"92"),
  1207 => (x"49",x"a2",x"c8",x"82"),
  1208 => (x"97",x"4b",x"a2",x"c9"),
  1209 => (x"97",x"1e",x"4b",x"6b"),
  1210 => (x"ca",x"1e",x"49",x"69"),
  1211 => (x"c0",x"49",x"12",x"82"),
  1212 => (x"c0",x"87",x"f0",x"f6"),
  1213 => (x"87",x"ce",x"d4",x"49"),
  1214 => (x"ca",x"c1",x"49",x"74"),
  1215 => (x"8e",x"f8",x"87",x"f9"),
  1216 => (x"1e",x"87",x"f8",x"f4"),
  1217 => (x"4b",x"71",x"1e",x"73"),
  1218 => (x"87",x"c3",x"ff",x"49"),
  1219 => (x"fe",x"fe",x"49",x"73"),
  1220 => (x"c1",x"49",x"c0",x"87"),
  1221 => (x"f4",x"87",x"c5",x"cc"),
  1222 => (x"73",x"1e",x"87",x"e3"),
  1223 => (x"c6",x"4b",x"71",x"1e"),
  1224 => (x"db",x"02",x"4a",x"a3"),
  1225 => (x"02",x"8a",x"c1",x"87"),
  1226 => (x"02",x"8a",x"87",x"d6"),
  1227 => (x"8a",x"87",x"da",x"c1"),
  1228 => (x"87",x"fc",x"c0",x"02"),
  1229 => (x"e1",x"c0",x"02",x"8a"),
  1230 => (x"cb",x"02",x"8a",x"87"),
  1231 => (x"87",x"db",x"c1",x"87"),
  1232 => (x"fa",x"fc",x"49",x"c7"),
  1233 => (x"87",x"de",x"c1",x"87"),
  1234 => (x"bf",x"c0",x"c1",x"c3"),
  1235 => (x"87",x"cb",x"c1",x"02"),
  1236 => (x"c3",x"88",x"c1",x"48"),
  1237 => (x"c1",x"58",x"c4",x"c1"),
  1238 => (x"c1",x"c3",x"87",x"c1"),
  1239 => (x"c0",x"02",x"bf",x"c4"),
  1240 => (x"c1",x"c3",x"87",x"f9"),
  1241 => (x"c1",x"48",x"bf",x"c0"),
  1242 => (x"c4",x"c1",x"c3",x"80"),
  1243 => (x"87",x"eb",x"c0",x"58"),
  1244 => (x"bf",x"c0",x"c1",x"c3"),
  1245 => (x"c3",x"89",x"c6",x"49"),
  1246 => (x"c0",x"59",x"c4",x"c1"),
  1247 => (x"da",x"03",x"a9",x"b7"),
  1248 => (x"c0",x"c1",x"c3",x"87"),
  1249 => (x"d2",x"78",x"c0",x"48"),
  1250 => (x"c4",x"c1",x"c3",x"87"),
  1251 => (x"87",x"cb",x"02",x"bf"),
  1252 => (x"bf",x"c0",x"c1",x"c3"),
  1253 => (x"c3",x"80",x"c6",x"48"),
  1254 => (x"c0",x"58",x"c4",x"c1"),
  1255 => (x"87",x"e6",x"d1",x"49"),
  1256 => (x"c8",x"c1",x"49",x"73"),
  1257 => (x"d4",x"f2",x"87",x"d1"),
  1258 => (x"5b",x"5e",x"0e",x"87"),
  1259 => (x"4c",x"71",x"0e",x"5c"),
  1260 => (x"74",x"1e",x"66",x"cc"),
  1261 => (x"c1",x"93",x"cb",x"4b"),
  1262 => (x"c4",x"83",x"f5",x"e3"),
  1263 => (x"49",x"6a",x"4a",x"a3"),
  1264 => (x"87",x"f4",x"f3",x"fe"),
  1265 => (x"7b",x"fd",x"c8",x"c1"),
  1266 => (x"d4",x"49",x"a3",x"c8"),
  1267 => (x"a3",x"c9",x"51",x"66"),
  1268 => (x"51",x"66",x"d8",x"49"),
  1269 => (x"dc",x"49",x"a3",x"ca"),
  1270 => (x"f1",x"26",x"51",x"66"),
  1271 => (x"5e",x"0e",x"87",x"dd"),
  1272 => (x"0e",x"5d",x"5c",x"5b"),
  1273 => (x"d8",x"86",x"d0",x"ff"),
  1274 => (x"a6",x"c4",x"59",x"a6"),
  1275 => (x"c4",x"78",x"c0",x"48"),
  1276 => (x"66",x"c4",x"c1",x"80"),
  1277 => (x"c1",x"80",x"c4",x"78"),
  1278 => (x"c1",x"80",x"c4",x"78"),
  1279 => (x"c4",x"c1",x"c3",x"78"),
  1280 => (x"c3",x"78",x"c1",x"48"),
  1281 => (x"48",x"bf",x"fc",x"c0"),
  1282 => (x"cb",x"05",x"a8",x"de"),
  1283 => (x"87",x"df",x"f3",x"87"),
  1284 => (x"a6",x"c8",x"49",x"70"),
  1285 => (x"87",x"f7",x"ce",x"59"),
  1286 => (x"e8",x"87",x"d6",x"e8"),
  1287 => (x"c5",x"e8",x"87",x"f8"),
  1288 => (x"c0",x"4c",x"70",x"87"),
  1289 => (x"c1",x"02",x"ac",x"fb"),
  1290 => (x"66",x"d4",x"87",x"d0"),
  1291 => (x"87",x"c2",x"c1",x"05"),
  1292 => (x"c1",x"1e",x"1e",x"c0"),
  1293 => (x"e8",x"e5",x"c1",x"1e"),
  1294 => (x"fd",x"49",x"c0",x"1e"),
  1295 => (x"d0",x"c1",x"87",x"eb"),
  1296 => (x"82",x"c4",x"4a",x"66"),
  1297 => (x"81",x"c7",x"49",x"6a"),
  1298 => (x"1e",x"c1",x"51",x"74"),
  1299 => (x"49",x"6a",x"1e",x"d8"),
  1300 => (x"d5",x"e8",x"81",x"c8"),
  1301 => (x"c1",x"86",x"d8",x"87"),
  1302 => (x"c0",x"48",x"66",x"c4"),
  1303 => (x"87",x"c7",x"01",x"a8"),
  1304 => (x"c1",x"48",x"a6",x"c4"),
  1305 => (x"c1",x"87",x"ce",x"78"),
  1306 => (x"c1",x"48",x"66",x"c4"),
  1307 => (x"58",x"a6",x"cc",x"88"),
  1308 => (x"e1",x"e7",x"87",x"c3"),
  1309 => (x"48",x"a6",x"cc",x"87"),
  1310 => (x"9c",x"74",x"78",x"c2"),
  1311 => (x"87",x"cb",x"cd",x"02"),
  1312 => (x"c1",x"48",x"66",x"c4"),
  1313 => (x"03",x"a8",x"66",x"c8"),
  1314 => (x"d8",x"87",x"c0",x"cd"),
  1315 => (x"78",x"c0",x"48",x"a6"),
  1316 => (x"70",x"87",x"d3",x"e6"),
  1317 => (x"ac",x"d0",x"c1",x"4c"),
  1318 => (x"87",x"d6",x"c2",x"05"),
  1319 => (x"e8",x"7e",x"66",x"d8"),
  1320 => (x"49",x"70",x"87",x"f7"),
  1321 => (x"e5",x"59",x"a6",x"dc"),
  1322 => (x"4c",x"70",x"87",x"fc"),
  1323 => (x"05",x"ac",x"ec",x"c0"),
  1324 => (x"c4",x"87",x"ea",x"c1"),
  1325 => (x"91",x"cb",x"49",x"66"),
  1326 => (x"81",x"66",x"c0",x"c1"),
  1327 => (x"6a",x"4a",x"a1",x"c4"),
  1328 => (x"4a",x"a1",x"c8",x"4d"),
  1329 => (x"c1",x"52",x"66",x"d8"),
  1330 => (x"e5",x"79",x"ff",x"c9"),
  1331 => (x"4c",x"70",x"87",x"d8"),
  1332 => (x"87",x"d8",x"02",x"9c"),
  1333 => (x"02",x"ac",x"fb",x"c0"),
  1334 => (x"55",x"74",x"87",x"d2"),
  1335 => (x"70",x"87",x"c7",x"e5"),
  1336 => (x"c7",x"02",x"9c",x"4c"),
  1337 => (x"ac",x"fb",x"c0",x"87"),
  1338 => (x"87",x"ee",x"ff",x"05"),
  1339 => (x"c2",x"55",x"e0",x"c0"),
  1340 => (x"97",x"c0",x"55",x"c1"),
  1341 => (x"49",x"66",x"d4",x"7d"),
  1342 => (x"db",x"05",x"a9",x"6e"),
  1343 => (x"48",x"66",x"c4",x"87"),
  1344 => (x"04",x"a8",x"66",x"c8"),
  1345 => (x"66",x"c4",x"87",x"ca"),
  1346 => (x"c8",x"80",x"c1",x"48"),
  1347 => (x"87",x"c8",x"58",x"a6"),
  1348 => (x"c1",x"48",x"66",x"c8"),
  1349 => (x"58",x"a6",x"cc",x"88"),
  1350 => (x"70",x"87",x"cb",x"e4"),
  1351 => (x"ac",x"d0",x"c1",x"4c"),
  1352 => (x"d0",x"87",x"c8",x"05"),
  1353 => (x"80",x"c1",x"48",x"66"),
  1354 => (x"c1",x"58",x"a6",x"d4"),
  1355 => (x"fd",x"02",x"ac",x"d0"),
  1356 => (x"a6",x"dc",x"87",x"ea"),
  1357 => (x"78",x"66",x"d4",x"48"),
  1358 => (x"dc",x"48",x"66",x"d8"),
  1359 => (x"c9",x"05",x"a8",x"66"),
  1360 => (x"e0",x"c0",x"87",x"db"),
  1361 => (x"f0",x"c0",x"48",x"a6"),
  1362 => (x"cc",x"80",x"c4",x"78"),
  1363 => (x"80",x"c4",x"78",x"66"),
  1364 => (x"74",x"7e",x"78",x"c0"),
  1365 => (x"88",x"fb",x"c0",x"48"),
  1366 => (x"58",x"a6",x"f0",x"c0"),
  1367 => (x"c8",x"02",x"98",x"70"),
  1368 => (x"cb",x"48",x"87",x"d6"),
  1369 => (x"a6",x"f0",x"c0",x"88"),
  1370 => (x"02",x"98",x"70",x"58"),
  1371 => (x"48",x"87",x"e9",x"c0"),
  1372 => (x"f0",x"c0",x"88",x"c9"),
  1373 => (x"98",x"70",x"58",x"a6"),
  1374 => (x"87",x"e1",x"c3",x"02"),
  1375 => (x"c0",x"88",x"c4",x"48"),
  1376 => (x"70",x"58",x"a6",x"f0"),
  1377 => (x"87",x"de",x"02",x"98"),
  1378 => (x"c0",x"88",x"c1",x"48"),
  1379 => (x"70",x"58",x"a6",x"f0"),
  1380 => (x"c8",x"c3",x"02",x"98"),
  1381 => (x"87",x"da",x"c7",x"87"),
  1382 => (x"48",x"a6",x"e0",x"c0"),
  1383 => (x"66",x"cc",x"78",x"c0"),
  1384 => (x"d0",x"80",x"c1",x"48"),
  1385 => (x"fd",x"e1",x"58",x"a6"),
  1386 => (x"c0",x"4c",x"70",x"87"),
  1387 => (x"d5",x"02",x"ac",x"ec"),
  1388 => (x"66",x"e0",x"c0",x"87"),
  1389 => (x"c0",x"87",x"c6",x"02"),
  1390 => (x"c9",x"5c",x"a6",x"e4"),
  1391 => (x"c0",x"48",x"74",x"87"),
  1392 => (x"e8",x"c0",x"88",x"f0"),
  1393 => (x"ec",x"c0",x"58",x"a6"),
  1394 => (x"87",x"cc",x"02",x"ac"),
  1395 => (x"70",x"87",x"d7",x"e1"),
  1396 => (x"ac",x"ec",x"c0",x"4c"),
  1397 => (x"87",x"f4",x"ff",x"05"),
  1398 => (x"1e",x"66",x"e0",x"c0"),
  1399 => (x"1e",x"49",x"66",x"d4"),
  1400 => (x"1e",x"66",x"ec",x"c0"),
  1401 => (x"1e",x"e8",x"e5",x"c1"),
  1402 => (x"f6",x"49",x"66",x"d4"),
  1403 => (x"1e",x"c0",x"87",x"fb"),
  1404 => (x"66",x"dc",x"1e",x"ca"),
  1405 => (x"c1",x"91",x"cb",x"49"),
  1406 => (x"d8",x"81",x"66",x"d8"),
  1407 => (x"a1",x"c4",x"48",x"a6"),
  1408 => (x"bf",x"66",x"d8",x"78"),
  1409 => (x"87",x"e2",x"e1",x"49"),
  1410 => (x"b7",x"c0",x"86",x"d8"),
  1411 => (x"c7",x"c1",x"06",x"a8"),
  1412 => (x"de",x"1e",x"c1",x"87"),
  1413 => (x"bf",x"66",x"c8",x"1e"),
  1414 => (x"87",x"ce",x"e1",x"49"),
  1415 => (x"49",x"70",x"86",x"c8"),
  1416 => (x"88",x"08",x"c0",x"48"),
  1417 => (x"58",x"a6",x"e4",x"c0"),
  1418 => (x"06",x"a8",x"b7",x"c0"),
  1419 => (x"c0",x"87",x"e9",x"c0"),
  1420 => (x"dd",x"48",x"66",x"e0"),
  1421 => (x"df",x"03",x"a8",x"b7"),
  1422 => (x"49",x"bf",x"6e",x"87"),
  1423 => (x"81",x"66",x"e0",x"c0"),
  1424 => (x"66",x"51",x"e0",x"c0"),
  1425 => (x"6e",x"81",x"c1",x"49"),
  1426 => (x"c1",x"c2",x"81",x"bf"),
  1427 => (x"66",x"e0",x"c0",x"51"),
  1428 => (x"6e",x"81",x"c2",x"49"),
  1429 => (x"51",x"c0",x"81",x"bf"),
  1430 => (x"db",x"c4",x"7e",x"c1"),
  1431 => (x"87",x"f9",x"e1",x"87"),
  1432 => (x"58",x"a6",x"e4",x"c0"),
  1433 => (x"c0",x"87",x"f2",x"e1"),
  1434 => (x"c0",x"58",x"a6",x"e8"),
  1435 => (x"c0",x"05",x"a8",x"ec"),
  1436 => (x"e4",x"c0",x"87",x"cb"),
  1437 => (x"e0",x"c0",x"48",x"a6"),
  1438 => (x"c4",x"c0",x"78",x"66"),
  1439 => (x"e5",x"de",x"ff",x"87"),
  1440 => (x"49",x"66",x"c4",x"87"),
  1441 => (x"c0",x"c1",x"91",x"cb"),
  1442 => (x"80",x"71",x"48",x"66"),
  1443 => (x"49",x"6e",x"7e",x"70"),
  1444 => (x"4a",x"6e",x"81",x"c8"),
  1445 => (x"e0",x"c0",x"82",x"ca"),
  1446 => (x"e4",x"c0",x"52",x"66"),
  1447 => (x"82",x"c1",x"4a",x"66"),
  1448 => (x"8a",x"66",x"e0",x"c0"),
  1449 => (x"30",x"72",x"48",x"c1"),
  1450 => (x"8a",x"c1",x"4a",x"70"),
  1451 => (x"97",x"79",x"97",x"72"),
  1452 => (x"c0",x"1e",x"49",x"69"),
  1453 => (x"c0",x"49",x"66",x"e4"),
  1454 => (x"c4",x"87",x"ea",x"e6"),
  1455 => (x"a6",x"f0",x"c0",x"86"),
  1456 => (x"c4",x"49",x"6e",x"58"),
  1457 => (x"dc",x"4d",x"69",x"81"),
  1458 => (x"66",x"d8",x"48",x"66"),
  1459 => (x"c8",x"c0",x"02",x"a8"),
  1460 => (x"48",x"a6",x"d8",x"87"),
  1461 => (x"c5",x"c0",x"78",x"c0"),
  1462 => (x"48",x"a6",x"d8",x"87"),
  1463 => (x"66",x"d8",x"78",x"c1"),
  1464 => (x"1e",x"e0",x"c0",x"1e"),
  1465 => (x"de",x"ff",x"49",x"75"),
  1466 => (x"86",x"c8",x"87",x"c0"),
  1467 => (x"b7",x"c0",x"4c",x"70"),
  1468 => (x"d4",x"c1",x"06",x"ac"),
  1469 => (x"c0",x"85",x"74",x"87"),
  1470 => (x"89",x"74",x"49",x"e0"),
  1471 => (x"e0",x"c1",x"4b",x"75"),
  1472 => (x"fe",x"71",x"4a",x"c3"),
  1473 => (x"c2",x"87",x"e1",x"e6"),
  1474 => (x"66",x"e8",x"c0",x"85"),
  1475 => (x"c0",x"80",x"c1",x"48"),
  1476 => (x"c0",x"58",x"a6",x"ec"),
  1477 => (x"c1",x"49",x"66",x"ec"),
  1478 => (x"02",x"a9",x"70",x"81"),
  1479 => (x"d8",x"87",x"c8",x"c0"),
  1480 => (x"78",x"c0",x"48",x"a6"),
  1481 => (x"d8",x"87",x"c5",x"c0"),
  1482 => (x"78",x"c1",x"48",x"a6"),
  1483 => (x"c2",x"1e",x"66",x"d8"),
  1484 => (x"e0",x"c0",x"49",x"a4"),
  1485 => (x"70",x"88",x"71",x"48"),
  1486 => (x"49",x"75",x"1e",x"49"),
  1487 => (x"87",x"ea",x"dc",x"ff"),
  1488 => (x"b7",x"c0",x"86",x"c8"),
  1489 => (x"c0",x"ff",x"01",x"a8"),
  1490 => (x"66",x"e8",x"c0",x"87"),
  1491 => (x"87",x"d1",x"c0",x"02"),
  1492 => (x"81",x"c9",x"49",x"6e"),
  1493 => (x"51",x"66",x"e8",x"c0"),
  1494 => (x"cb",x"c1",x"48",x"6e"),
  1495 => (x"cc",x"c0",x"78",x"cf"),
  1496 => (x"c9",x"49",x"6e",x"87"),
  1497 => (x"6e",x"51",x"c2",x"81"),
  1498 => (x"c3",x"cc",x"c1",x"48"),
  1499 => (x"c0",x"7e",x"c1",x"78"),
  1500 => (x"db",x"ff",x"87",x"c6"),
  1501 => (x"4c",x"70",x"87",x"e0"),
  1502 => (x"f5",x"c0",x"02",x"6e"),
  1503 => (x"48",x"66",x"c4",x"87"),
  1504 => (x"04",x"a8",x"66",x"c8"),
  1505 => (x"c4",x"87",x"cb",x"c0"),
  1506 => (x"80",x"c1",x"48",x"66"),
  1507 => (x"c0",x"58",x"a6",x"c8"),
  1508 => (x"66",x"c8",x"87",x"e0"),
  1509 => (x"cc",x"88",x"c1",x"48"),
  1510 => (x"d5",x"c0",x"58",x"a6"),
  1511 => (x"ac",x"c6",x"c1",x"87"),
  1512 => (x"87",x"c8",x"c0",x"05"),
  1513 => (x"c1",x"48",x"66",x"cc"),
  1514 => (x"58",x"a6",x"d0",x"80"),
  1515 => (x"87",x"e6",x"da",x"ff"),
  1516 => (x"66",x"d0",x"4c",x"70"),
  1517 => (x"d4",x"80",x"c1",x"48"),
  1518 => (x"9c",x"74",x"58",x"a6"),
  1519 => (x"87",x"cb",x"c0",x"02"),
  1520 => (x"c1",x"48",x"66",x"c4"),
  1521 => (x"04",x"a8",x"66",x"c8"),
  1522 => (x"ff",x"87",x"c0",x"f3"),
  1523 => (x"c4",x"87",x"fe",x"d9"),
  1524 => (x"a8",x"c7",x"48",x"66"),
  1525 => (x"87",x"e5",x"c0",x"03"),
  1526 => (x"48",x"c4",x"c1",x"c3"),
  1527 => (x"66",x"c4",x"78",x"c0"),
  1528 => (x"c1",x"91",x"cb",x"49"),
  1529 => (x"c4",x"81",x"66",x"c0"),
  1530 => (x"4a",x"6a",x"4a",x"a1"),
  1531 => (x"c4",x"79",x"52",x"c0"),
  1532 => (x"80",x"c1",x"48",x"66"),
  1533 => (x"c7",x"58",x"a6",x"c8"),
  1534 => (x"db",x"ff",x"04",x"a8"),
  1535 => (x"8e",x"d0",x"ff",x"87"),
  1536 => (x"3a",x"87",x"f6",x"e0"),
  1537 => (x"73",x"1e",x"00",x"20"),
  1538 => (x"9b",x"4b",x"71",x"1e"),
  1539 => (x"c3",x"87",x"c6",x"02"),
  1540 => (x"c0",x"48",x"c0",x"c1"),
  1541 => (x"c3",x"1e",x"c7",x"78"),
  1542 => (x"49",x"bf",x"c0",x"c1"),
  1543 => (x"f5",x"e3",x"c1",x"1e"),
  1544 => (x"fc",x"c0",x"c3",x"1e"),
  1545 => (x"f5",x"ee",x"49",x"bf"),
  1546 => (x"c3",x"86",x"cc",x"87"),
  1547 => (x"49",x"bf",x"fc",x"c0"),
  1548 => (x"73",x"87",x"f4",x"e9"),
  1549 => (x"87",x"c8",x"02",x"9b"),
  1550 => (x"49",x"f5",x"e3",x"c1"),
  1551 => (x"87",x"c9",x"f7",x"c0"),
  1552 => (x"87",x"f9",x"df",x"ff"),
  1553 => (x"f3",x"f2",x"c2",x"1e"),
  1554 => (x"c1",x"50",x"c0",x"48"),
  1555 => (x"49",x"bf",x"d8",x"e5"),
  1556 => (x"87",x"f4",x"cc",x"c1"),
  1557 => (x"4f",x"26",x"48",x"c0"),
  1558 => (x"87",x"df",x"cd",x"1e"),
  1559 => (x"e5",x"fe",x"49",x"c1"),
  1560 => (x"d6",x"e9",x"fe",x"87"),
  1561 => (x"02",x"98",x"70",x"87"),
  1562 => (x"f2",x"fe",x"87",x"cd"),
  1563 => (x"98",x"70",x"87",x"d3"),
  1564 => (x"c1",x"87",x"c4",x"02"),
  1565 => (x"c0",x"87",x"c2",x"4a"),
  1566 => (x"05",x"9a",x"72",x"4a"),
  1567 => (x"1e",x"c0",x"87",x"ce"),
  1568 => (x"49",x"e8",x"e2",x"c1"),
  1569 => (x"87",x"de",x"c2",x"c1"),
  1570 => (x"87",x"fe",x"86",x"c4"),
  1571 => (x"e2",x"c1",x"1e",x"c0"),
  1572 => (x"c2",x"c1",x"49",x"f3"),
  1573 => (x"1e",x"c0",x"87",x"d0"),
  1574 => (x"70",x"87",x"e9",x"fe"),
  1575 => (x"c5",x"c2",x"c1",x"49"),
  1576 => (x"87",x"e2",x"c3",x"87"),
  1577 => (x"4f",x"26",x"8e",x"f8"),
  1578 => (x"66",x"20",x"44",x"53"),
  1579 => (x"65",x"6c",x"69",x"61"),
  1580 => (x"42",x"00",x"2e",x"64"),
  1581 => (x"69",x"74",x"6f",x"6f"),
  1582 => (x"2e",x"2e",x"67",x"6e"),
  1583 => (x"c0",x"1e",x"00",x"2e"),
  1584 => (x"87",x"ce",x"d5",x"49"),
  1585 => (x"87",x"e1",x"f9",x"c0"),
  1586 => (x"87",x"d0",x"c5",x"c1"),
  1587 => (x"4f",x"26",x"87",x"f1"),
  1588 => (x"c0",x"c1",x"c3",x"1e"),
  1589 => (x"c3",x"78",x"c0",x"48"),
  1590 => (x"c0",x"48",x"fc",x"c0"),
  1591 => (x"87",x"f8",x"fd",x"78"),
  1592 => (x"c0",x"87",x"db",x"ff"),
  1593 => (x"80",x"4f",x"26",x"48"),
  1594 => (x"69",x"78",x"45",x"20"),
  1595 => (x"20",x"80",x"00",x"74"),
  1596 => (x"6b",x"63",x"61",x"42"),
  1597 => (x"00",x"12",x"7f",x"00"),
  1598 => (x"00",x"30",x"55",x"00"),
  1599 => (x"00",x"00",x"00",x"00"),
  1600 => (x"00",x"00",x"12",x"7f"),
  1601 => (x"00",x"00",x"30",x"73"),
  1602 => (x"7f",x"00",x"00",x"00"),
  1603 => (x"91",x"00",x"00",x"12"),
  1604 => (x"00",x"00",x"00",x"30"),
  1605 => (x"12",x"7f",x"00",x"00"),
  1606 => (x"30",x"af",x"00",x"00"),
  1607 => (x"00",x"00",x"00",x"00"),
  1608 => (x"00",x"12",x"7f",x"00"),
  1609 => (x"00",x"30",x"cd",x"00"),
  1610 => (x"00",x"00",x"00",x"00"),
  1611 => (x"00",x"00",x"12",x"7f"),
  1612 => (x"00",x"00",x"30",x"eb"),
  1613 => (x"7f",x"00",x"00",x"00"),
  1614 => (x"09",x"00",x"00",x"12"),
  1615 => (x"00",x"00",x"00",x"31"),
  1616 => (x"12",x"7f",x"00",x"00"),
  1617 => (x"00",x"00",x"00",x"00"),
  1618 => (x"00",x"00",x"00",x"00"),
  1619 => (x"00",x"13",x"1a",x"00"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"00",x"00",x"00",x"00"),
  1622 => (x"00",x"00",x"19",x"5c"),
  1623 => (x"54",x"4f",x"4f",x"42"),
  1624 => (x"20",x"20",x"20",x"20"),
  1625 => (x"00",x"4d",x"4f",x"52"),
  1626 => (x"64",x"61",x"6f",x"4c"),
  1627 => (x"00",x"2e",x"2a",x"20"),
  1628 => (x"48",x"f0",x"fe",x"1e"),
  1629 => (x"09",x"cd",x"78",x"c0"),
  1630 => (x"4f",x"26",x"09",x"79"),
  1631 => (x"f0",x"fe",x"1e",x"1e"),
  1632 => (x"26",x"48",x"7e",x"bf"),
  1633 => (x"fe",x"1e",x"4f",x"26"),
  1634 => (x"78",x"c1",x"48",x"f0"),
  1635 => (x"fe",x"1e",x"4f",x"26"),
  1636 => (x"78",x"c0",x"48",x"f0"),
  1637 => (x"71",x"1e",x"4f",x"26"),
  1638 => (x"7a",x"97",x"c0",x"4a"),
  1639 => (x"c0",x"49",x"a2",x"c1"),
  1640 => (x"49",x"a2",x"ca",x"51"),
  1641 => (x"a2",x"cb",x"51",x"c0"),
  1642 => (x"26",x"51",x"c0",x"49"),
  1643 => (x"5b",x"5e",x"0e",x"4f"),
  1644 => (x"86",x"f0",x"0e",x"5c"),
  1645 => (x"a4",x"ca",x"4c",x"71"),
  1646 => (x"7e",x"69",x"97",x"49"),
  1647 => (x"97",x"4b",x"a4",x"cb"),
  1648 => (x"a6",x"c8",x"48",x"6b"),
  1649 => (x"cc",x"80",x"c1",x"58"),
  1650 => (x"98",x"c7",x"58",x"a6"),
  1651 => (x"6e",x"58",x"a6",x"d0"),
  1652 => (x"a8",x"66",x"cc",x"48"),
  1653 => (x"97",x"87",x"db",x"05"),
  1654 => (x"6b",x"97",x"7e",x"69"),
  1655 => (x"58",x"a6",x"c8",x"48"),
  1656 => (x"a6",x"cc",x"80",x"c1"),
  1657 => (x"d0",x"98",x"c7",x"58"),
  1658 => (x"48",x"6e",x"58",x"a6"),
  1659 => (x"02",x"a8",x"66",x"cc"),
  1660 => (x"d9",x"fe",x"87",x"e5"),
  1661 => (x"4a",x"a4",x"cc",x"87"),
  1662 => (x"72",x"49",x"6b",x"97"),
  1663 => (x"66",x"dc",x"49",x"a1"),
  1664 => (x"7e",x"6b",x"97",x"51"),
  1665 => (x"80",x"c1",x"48",x"6e"),
  1666 => (x"c7",x"58",x"a6",x"c8"),
  1667 => (x"58",x"a6",x"cc",x"98"),
  1668 => (x"c3",x"7b",x"97",x"70"),
  1669 => (x"ed",x"fd",x"87",x"d2"),
  1670 => (x"c2",x"8e",x"f0",x"87"),
  1671 => (x"26",x"4d",x"26",x"87"),
  1672 => (x"26",x"4b",x"26",x"4c"),
  1673 => (x"5b",x"5e",x"0e",x"4f"),
  1674 => (x"f4",x"0e",x"5d",x"5c"),
  1675 => (x"97",x"4d",x"71",x"86"),
  1676 => (x"a5",x"c1",x"7e",x"6d"),
  1677 => (x"48",x"6c",x"97",x"4c"),
  1678 => (x"6e",x"58",x"a6",x"c8"),
  1679 => (x"a8",x"66",x"c4",x"48"),
  1680 => (x"ff",x"87",x"c5",x"05"),
  1681 => (x"87",x"e6",x"c0",x"48"),
  1682 => (x"c2",x"87",x"c3",x"fd"),
  1683 => (x"6c",x"97",x"49",x"a5"),
  1684 => (x"4b",x"a3",x"71",x"4b"),
  1685 => (x"97",x"4b",x"6b",x"97"),
  1686 => (x"48",x"6e",x"7e",x"6c"),
  1687 => (x"a6",x"c8",x"80",x"c1"),
  1688 => (x"cc",x"98",x"c7",x"58"),
  1689 => (x"97",x"70",x"58",x"a6"),
  1690 => (x"87",x"da",x"fc",x"7c"),
  1691 => (x"8e",x"f4",x"48",x"73"),
  1692 => (x"0e",x"87",x"ea",x"fe"),
  1693 => (x"0e",x"5c",x"5b",x"5e"),
  1694 => (x"4c",x"71",x"86",x"f4"),
  1695 => (x"c3",x"4a",x"66",x"d8"),
  1696 => (x"a4",x"c2",x"9a",x"ff"),
  1697 => (x"49",x"6c",x"97",x"4b"),
  1698 => (x"72",x"49",x"a1",x"73"),
  1699 => (x"7e",x"6c",x"97",x"51"),
  1700 => (x"80",x"c1",x"48",x"6e"),
  1701 => (x"c7",x"58",x"a6",x"c8"),
  1702 => (x"58",x"a6",x"cc",x"98"),
  1703 => (x"8e",x"f4",x"54",x"70"),
  1704 => (x"1e",x"87",x"fc",x"fd"),
  1705 => (x"69",x"97",x"86",x"f0"),
  1706 => (x"4a",x"a1",x"c1",x"7e"),
  1707 => (x"c8",x"48",x"6a",x"97"),
  1708 => (x"48",x"6e",x"58",x"a6"),
  1709 => (x"a8",x"b7",x"66",x"c4"),
  1710 => (x"97",x"87",x"d3",x"04"),
  1711 => (x"6a",x"97",x"7e",x"69"),
  1712 => (x"58",x"a6",x"c8",x"48"),
  1713 => (x"66",x"c4",x"48",x"6e"),
  1714 => (x"58",x"a6",x"cc",x"88"),
  1715 => (x"7e",x"11",x"87",x"d6"),
  1716 => (x"80",x"c8",x"48",x"6e"),
  1717 => (x"48",x"12",x"58",x"a6"),
  1718 => (x"c4",x"58",x"a6",x"cc"),
  1719 => (x"66",x"c8",x"48",x"66"),
  1720 => (x"58",x"a6",x"d0",x"88"),
  1721 => (x"4f",x"26",x"8e",x"f0"),
  1722 => (x"f4",x"1e",x"73",x"1e"),
  1723 => (x"87",x"de",x"fa",x"86"),
  1724 => (x"49",x"4b",x"bf",x"e0"),
  1725 => (x"99",x"c0",x"e0",x"c0"),
  1726 => (x"73",x"87",x"cb",x"02"),
  1727 => (x"e7",x"c4",x"c3",x"1e"),
  1728 => (x"87",x"ef",x"fd",x"49"),
  1729 => (x"49",x"73",x"86",x"c4"),
  1730 => (x"02",x"99",x"c0",x"d0"),
  1731 => (x"c3",x"87",x"c0",x"c1"),
  1732 => (x"bf",x"97",x"f1",x"c4"),
  1733 => (x"f2",x"c4",x"c3",x"7e"),
  1734 => (x"c8",x"48",x"bf",x"97"),
  1735 => (x"48",x"6e",x"58",x"a6"),
  1736 => (x"02",x"a8",x"66",x"c4"),
  1737 => (x"c3",x"87",x"e8",x"c0"),
  1738 => (x"bf",x"97",x"f1",x"c4"),
  1739 => (x"f3",x"c4",x"c3",x"49"),
  1740 => (x"e0",x"48",x"11",x"81"),
  1741 => (x"c4",x"c3",x"78",x"08"),
  1742 => (x"7e",x"bf",x"97",x"f1"),
  1743 => (x"80",x"c1",x"48",x"6e"),
  1744 => (x"c7",x"58",x"a6",x"c8"),
  1745 => (x"58",x"a6",x"cc",x"98"),
  1746 => (x"48",x"f1",x"c4",x"c3"),
  1747 => (x"e4",x"50",x"66",x"c8"),
  1748 => (x"c0",x"49",x"4b",x"bf"),
  1749 => (x"02",x"99",x"c0",x"e0"),
  1750 => (x"1e",x"73",x"87",x"cb"),
  1751 => (x"49",x"fb",x"c4",x"c3"),
  1752 => (x"c4",x"87",x"d0",x"fc"),
  1753 => (x"d0",x"49",x"73",x"86"),
  1754 => (x"c1",x"02",x"99",x"c0"),
  1755 => (x"c5",x"c3",x"87",x"c0"),
  1756 => (x"7e",x"bf",x"97",x"c5"),
  1757 => (x"97",x"c6",x"c5",x"c3"),
  1758 => (x"a6",x"c8",x"48",x"bf"),
  1759 => (x"c4",x"48",x"6e",x"58"),
  1760 => (x"c0",x"02",x"a8",x"66"),
  1761 => (x"c5",x"c3",x"87",x"e8"),
  1762 => (x"49",x"bf",x"97",x"c5"),
  1763 => (x"81",x"c7",x"c5",x"c3"),
  1764 => (x"08",x"e4",x"48",x"11"),
  1765 => (x"c5",x"c5",x"c3",x"78"),
  1766 => (x"6e",x"7e",x"bf",x"97"),
  1767 => (x"c8",x"80",x"c1",x"48"),
  1768 => (x"98",x"c7",x"58",x"a6"),
  1769 => (x"c3",x"58",x"a6",x"cc"),
  1770 => (x"c8",x"48",x"c5",x"c5"),
  1771 => (x"cb",x"f7",x"50",x"66"),
  1772 => (x"f7",x"7e",x"70",x"87"),
  1773 => (x"8e",x"f4",x"87",x"d0"),
  1774 => (x"1e",x"87",x"e6",x"f9"),
  1775 => (x"49",x"e7",x"c4",x"c3"),
  1776 => (x"c3",x"87",x"d3",x"f7"),
  1777 => (x"f7",x"49",x"fb",x"c4"),
  1778 => (x"eb",x"c1",x"87",x"cc"),
  1779 => (x"df",x"f6",x"49",x"e8"),
  1780 => (x"87",x"d9",x"c5",x"87"),
  1781 => (x"5e",x"0e",x"4f",x"26"),
  1782 => (x"0e",x"5d",x"5c",x"5b"),
  1783 => (x"bf",x"ec",x"c5",x"c3"),
  1784 => (x"ea",x"f0",x"c1",x"4a"),
  1785 => (x"72",x"4c",x"49",x"bf"),
  1786 => (x"f6",x"4d",x"71",x"bc"),
  1787 => (x"4b",x"c0",x"87",x"e0"),
  1788 => (x"99",x"d0",x"49",x"74"),
  1789 => (x"75",x"87",x"d5",x"02"),
  1790 => (x"71",x"99",x"d0",x"49"),
  1791 => (x"c1",x"1e",x"c0",x"1e"),
  1792 => (x"73",x"4a",x"fc",x"f6"),
  1793 => (x"c0",x"49",x"12",x"82"),
  1794 => (x"86",x"c8",x"87",x"e4"),
  1795 => (x"83",x"2d",x"2c",x"c1"),
  1796 => (x"ff",x"04",x"ab",x"c8"),
  1797 => (x"ed",x"f5",x"87",x"da"),
  1798 => (x"ea",x"f0",x"c1",x"87"),
  1799 => (x"ec",x"c5",x"c3",x"48"),
  1800 => (x"4d",x"26",x"78",x"bf"),
  1801 => (x"4b",x"26",x"4c",x"26"),
  1802 => (x"00",x"00",x"4f",x"26"),
  1803 => (x"ff",x"1e",x"00",x"00"),
  1804 => (x"e1",x"c8",x"48",x"d0"),
  1805 => (x"48",x"d4",x"ff",x"78"),
  1806 => (x"66",x"c4",x"78",x"c5"),
  1807 => (x"c3",x"87",x"c3",x"02"),
  1808 => (x"66",x"c8",x"78",x"e0"),
  1809 => (x"ff",x"87",x"c6",x"02"),
  1810 => (x"f0",x"c3",x"48",x"d4"),
  1811 => (x"48",x"d4",x"ff",x"78"),
  1812 => (x"d0",x"ff",x"78",x"71"),
  1813 => (x"78",x"e1",x"c8",x"48"),
  1814 => (x"26",x"78",x"e0",x"c0"),
  1815 => (x"5b",x"5e",x"0e",x"4f"),
  1816 => (x"4c",x"71",x"0e",x"5c"),
  1817 => (x"49",x"e7",x"c4",x"c3"),
  1818 => (x"70",x"87",x"fa",x"f6"),
  1819 => (x"aa",x"b7",x"c0",x"4a"),
  1820 => (x"87",x"e3",x"c2",x"04"),
  1821 => (x"05",x"aa",x"e0",x"c3"),
  1822 => (x"f4",x"c1",x"87",x"c9"),
  1823 => (x"78",x"c1",x"48",x"e0"),
  1824 => (x"c3",x"87",x"d4",x"c2"),
  1825 => (x"c9",x"05",x"aa",x"f0"),
  1826 => (x"dc",x"f4",x"c1",x"87"),
  1827 => (x"c1",x"78",x"c1",x"48"),
  1828 => (x"f4",x"c1",x"87",x"f5"),
  1829 => (x"c7",x"02",x"bf",x"e0"),
  1830 => (x"c2",x"4b",x"72",x"87"),
  1831 => (x"87",x"c2",x"b3",x"c0"),
  1832 => (x"9c",x"74",x"4b",x"72"),
  1833 => (x"c1",x"87",x"d1",x"05"),
  1834 => (x"1e",x"bf",x"dc",x"f4"),
  1835 => (x"bf",x"e0",x"f4",x"c1"),
  1836 => (x"fd",x"49",x"72",x"1e"),
  1837 => (x"86",x"c8",x"87",x"f8"),
  1838 => (x"bf",x"dc",x"f4",x"c1"),
  1839 => (x"87",x"e0",x"c0",x"02"),
  1840 => (x"b7",x"c4",x"49",x"73"),
  1841 => (x"f5",x"c1",x"91",x"29"),
  1842 => (x"4a",x"73",x"81",x"fc"),
  1843 => (x"92",x"c2",x"9a",x"cf"),
  1844 => (x"30",x"72",x"48",x"c1"),
  1845 => (x"ba",x"ff",x"4a",x"70"),
  1846 => (x"98",x"69",x"48",x"72"),
  1847 => (x"87",x"db",x"79",x"70"),
  1848 => (x"b7",x"c4",x"49",x"73"),
  1849 => (x"f5",x"c1",x"91",x"29"),
  1850 => (x"4a",x"73",x"81",x"fc"),
  1851 => (x"92",x"c2",x"9a",x"cf"),
  1852 => (x"30",x"72",x"48",x"c3"),
  1853 => (x"69",x"48",x"4a",x"70"),
  1854 => (x"c1",x"79",x"70",x"b0"),
  1855 => (x"c0",x"48",x"e0",x"f4"),
  1856 => (x"dc",x"f4",x"c1",x"78"),
  1857 => (x"c3",x"78",x"c0",x"48"),
  1858 => (x"f4",x"49",x"e7",x"c4"),
  1859 => (x"4a",x"70",x"87",x"d7"),
  1860 => (x"03",x"aa",x"b7",x"c0"),
  1861 => (x"c0",x"87",x"dd",x"fd"),
  1862 => (x"87",x"c8",x"fc",x"48"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"49",x"4a",x"71",x"1e"),
  1866 => (x"26",x"87",x"f2",x"fc"),
  1867 => (x"4a",x"c0",x"1e",x"4f"),
  1868 => (x"91",x"c4",x"49",x"72"),
  1869 => (x"81",x"fc",x"f5",x"c1"),
  1870 => (x"82",x"c1",x"79",x"c0"),
  1871 => (x"04",x"aa",x"b7",x"d0"),
  1872 => (x"4f",x"26",x"87",x"ee"),
  1873 => (x"5c",x"5b",x"5e",x"0e"),
  1874 => (x"4d",x"71",x"0e",x"5d"),
  1875 => (x"75",x"87",x"ff",x"f0"),
  1876 => (x"2a",x"b7",x"c4",x"4a"),
  1877 => (x"fc",x"f5",x"c1",x"92"),
  1878 => (x"cf",x"4c",x"75",x"82"),
  1879 => (x"6a",x"94",x"c2",x"9c"),
  1880 => (x"2b",x"74",x"4b",x"49"),
  1881 => (x"48",x"c2",x"9b",x"c3"),
  1882 => (x"4c",x"70",x"30",x"74"),
  1883 => (x"48",x"74",x"bc",x"ff"),
  1884 => (x"7a",x"70",x"98",x"71"),
  1885 => (x"73",x"87",x"cf",x"f0"),
  1886 => (x"87",x"e6",x"fa",x"48"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"00",x"00",x"00",x"00"),
  1894 => (x"00",x"00",x"00",x"00"),
  1895 => (x"00",x"00",x"00",x"00"),
  1896 => (x"00",x"00",x"00",x"00"),
  1897 => (x"00",x"00",x"00",x"00"),
  1898 => (x"00",x"00",x"00",x"00"),
  1899 => (x"00",x"00",x"00",x"00"),
  1900 => (x"00",x"00",x"00",x"00"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"25",x"26",x"1e",x"16"),
  1904 => (x"3e",x"3d",x"36",x"2e"),
  1905 => (x"71",x"1e",x"73",x"1e"),
  1906 => (x"fb",x"c4",x"c3",x"4b"),
  1907 => (x"87",x"d5",x"f1",x"49"),
  1908 => (x"c4",x"1e",x"49",x"70"),
  1909 => (x"87",x"c4",x"c8",x"49"),
  1910 => (x"c4",x"c3",x"86",x"c4"),
  1911 => (x"c4",x"f1",x"49",x"fb"),
  1912 => (x"ff",x"49",x"70",x"87"),
  1913 => (x"78",x"71",x"48",x"d4"),
  1914 => (x"49",x"fb",x"c4",x"c3"),
  1915 => (x"70",x"87",x"f6",x"f0"),
  1916 => (x"48",x"d4",x"ff",x"49"),
  1917 => (x"d0",x"ff",x"78",x"71"),
  1918 => (x"78",x"e0",x"c0",x"48"),
  1919 => (x"c7",x"05",x"ab",x"c4"),
  1920 => (x"fb",x"c4",x"c3",x"87"),
  1921 => (x"87",x"dd",x"f0",x"49"),
  1922 => (x"4d",x"26",x"87",x"c4"),
  1923 => (x"4b",x"26",x"4c",x"26"),
  1924 => (x"5e",x"0e",x"4f",x"26"),
  1925 => (x"0e",x"5d",x"5c",x"5b"),
  1926 => (x"02",x"9a",x"4a",x"71"),
  1927 => (x"fe",x"c1",x"87",x"c6"),
  1928 => (x"78",x"c0",x"48",x"ed"),
  1929 => (x"bf",x"ed",x"fe",x"c1"),
  1930 => (x"87",x"c6",x"c1",x"05"),
  1931 => (x"49",x"fb",x"c4",x"c3"),
  1932 => (x"c0",x"87",x"f2",x"ef"),
  1933 => (x"cd",x"04",x"a8",x"b7"),
  1934 => (x"fb",x"c4",x"c3",x"87"),
  1935 => (x"87",x"e5",x"ef",x"49"),
  1936 => (x"03",x"a8",x"b7",x"c0"),
  1937 => (x"fe",x"c1",x"87",x"f3"),
  1938 => (x"c1",x"49",x"bf",x"ed"),
  1939 => (x"c1",x"48",x"ed",x"fe"),
  1940 => (x"fe",x"c1",x"78",x"a1"),
  1941 => (x"48",x"11",x"81",x"fd"),
  1942 => (x"58",x"f5",x"fe",x"c1"),
  1943 => (x"48",x"f5",x"fe",x"c1"),
  1944 => (x"f2",x"c0",x"78",x"c0"),
  1945 => (x"da",x"ec",x"c0",x"49"),
  1946 => (x"c3",x"49",x"70",x"87"),
  1947 => (x"c4",x"59",x"d3",x"c5"),
  1948 => (x"fe",x"c1",x"87",x"f8"),
  1949 => (x"c1",x"02",x"bf",x"f5"),
  1950 => (x"c4",x"c3",x"87",x"f2"),
  1951 => (x"e4",x"ee",x"49",x"fb"),
  1952 => (x"a8",x"b7",x"c0",x"87"),
  1953 => (x"c1",x"87",x"cd",x"04"),
  1954 => (x"48",x"bf",x"f5",x"fe"),
  1955 => (x"fe",x"c1",x"88",x"c1"),
  1956 => (x"87",x"db",x"58",x"f9"),
  1957 => (x"bf",x"cf",x"c5",x"c3"),
  1958 => (x"f2",x"eb",x"c0",x"49"),
  1959 => (x"02",x"98",x"70",x"87"),
  1960 => (x"c4",x"c3",x"87",x"cd"),
  1961 => (x"ed",x"eb",x"49",x"fb"),
  1962 => (x"ed",x"fe",x"c1",x"87"),
  1963 => (x"c1",x"78",x"c0",x"48"),
  1964 => (x"05",x"bf",x"f1",x"fe"),
  1965 => (x"c1",x"87",x"f3",x"c3"),
  1966 => (x"05",x"bf",x"f5",x"fe"),
  1967 => (x"c1",x"87",x"eb",x"c3"),
  1968 => (x"49",x"bf",x"ed",x"fe"),
  1969 => (x"48",x"ed",x"fe",x"c1"),
  1970 => (x"c1",x"78",x"a1",x"c1"),
  1971 => (x"11",x"81",x"fd",x"fe"),
  1972 => (x"c0",x"c2",x"49",x"4b"),
  1973 => (x"cc",x"c0",x"02",x"99"),
  1974 => (x"c1",x"48",x"73",x"87"),
  1975 => (x"fe",x"c1",x"98",x"ff"),
  1976 => (x"c5",x"c3",x"58",x"f9"),
  1977 => (x"f5",x"fe",x"c1",x"87"),
  1978 => (x"87",x"fe",x"c2",x"5b"),
  1979 => (x"bf",x"f1",x"fe",x"c1"),
  1980 => (x"87",x"db",x"c1",x"02"),
  1981 => (x"bf",x"cf",x"c5",x"c3"),
  1982 => (x"d2",x"ea",x"c0",x"49"),
  1983 => (x"02",x"98",x"70",x"87"),
  1984 => (x"c1",x"87",x"e7",x"c2"),
  1985 => (x"49",x"bf",x"ed",x"fe"),
  1986 => (x"48",x"ed",x"fe",x"c1"),
  1987 => (x"c1",x"78",x"a1",x"c1"),
  1988 => (x"97",x"81",x"fd",x"fe"),
  1989 => (x"c3",x"1e",x"49",x"69"),
  1990 => (x"ea",x"49",x"fb",x"c4"),
  1991 => (x"86",x"c4",x"87",x"cf"),
  1992 => (x"bf",x"f1",x"fe",x"c1"),
  1993 => (x"c1",x"89",x"c1",x"49"),
  1994 => (x"c1",x"59",x"f5",x"fe"),
  1995 => (x"c1",x"48",x"f5",x"fe"),
  1996 => (x"02",x"99",x"71",x"78"),
  1997 => (x"c0",x"87",x"c6",x"c0"),
  1998 => (x"c3",x"c0",x"4c",x"f2"),
  1999 => (x"4c",x"dc",x"d7",x"87"),
  2000 => (x"e8",x"c0",x"49",x"74"),
  2001 => (x"49",x"70",x"87",x"fd"),
  2002 => (x"59",x"d3",x"c5",x"c3"),
  2003 => (x"c3",x"87",x"db",x"c1"),
  2004 => (x"ed",x"49",x"fb",x"c4"),
  2005 => (x"4b",x"70",x"87",x"cd"),
  2006 => (x"ee",x"c0",x"02",x"9b"),
  2007 => (x"f9",x"fe",x"c1",x"87"),
  2008 => (x"03",x"ab",x"b7",x"bf"),
  2009 => (x"c3",x"87",x"e4",x"c0"),
  2010 => (x"49",x"bf",x"cf",x"c5"),
  2011 => (x"87",x"df",x"e8",x"c0"),
  2012 => (x"c0",x"02",x"98",x"70"),
  2013 => (x"48",x"c7",x"87",x"f4"),
  2014 => (x"bf",x"f9",x"fe",x"c1"),
  2015 => (x"fd",x"fe",x"c1",x"88"),
  2016 => (x"fb",x"c4",x"c3",x"58"),
  2017 => (x"87",x"ce",x"e8",x"49"),
  2018 => (x"d7",x"87",x"df",x"c0"),
  2019 => (x"e7",x"c0",x"49",x"dc"),
  2020 => (x"49",x"70",x"87",x"f1"),
  2021 => (x"59",x"d3",x"c5",x"c3"),
  2022 => (x"bf",x"f9",x"fe",x"c1"),
  2023 => (x"04",x"ab",x"b7",x"4a"),
  2024 => (x"49",x"87",x"c7",x"c0"),
  2025 => (x"fe",x"87",x"dd",x"f8"),
  2026 => (x"dd",x"f9",x"87",x"e5"),
  2027 => (x"00",x"00",x"00",x"87"),
  2028 => (x"00",x"00",x"00",x"00"),
  2029 => (x"00",x"00",x"00",x"00"),
  2030 => (x"00",x"00",x"04",x"00"),
  2031 => (x"82",x"ff",x"01",x"00"),
  2032 => (x"f3",x"c8",x"f3",x"08"),
  2033 => (x"f2",x"50",x"f3",x"64"),
  2034 => (x"f4",x"01",x"81",x"01"),
  2035 => (x"d0",x"ff",x"1e",x"00"),
  2036 => (x"78",x"e1",x"c8",x"48"),
  2037 => (x"d4",x"ff",x"48",x"71"),
  2038 => (x"4f",x"26",x"78",x"08"),
  2039 => (x"48",x"d0",x"ff",x"1e"),
  2040 => (x"71",x"78",x"e1",x"c8"),
  2041 => (x"08",x"d4",x"ff",x"48"),
  2042 => (x"48",x"66",x"c4",x"78"),
  2043 => (x"78",x"08",x"d4",x"ff"),
  2044 => (x"71",x"1e",x"4f",x"26"),
  2045 => (x"49",x"66",x"c4",x"4a"),
  2046 => (x"ff",x"49",x"72",x"1e"),
  2047 => (x"d0",x"ff",x"87",x"de"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

