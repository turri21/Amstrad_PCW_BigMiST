library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e8c8c387",
    12 => x"86c0c64e",
    13 => x"49e8c8c3",
    14 => x"48e4f3c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c5e2",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfe4f3",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"f3c21e73",
   176 => x"78c148e4",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"e8f3c287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58ecf3c2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49ecf3",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"f3c287f8",
   280 => x"49bf97ec",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"f3c287e7",
   284 => x"49bf97f3",
   285 => x"f3c231d0",
   286 => x"4abf97f4",
   287 => x"b17232c8",
   288 => x"97f5f3c2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"f5f3c287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97f6f3",
   297 => x"2ab7c74a",
   298 => x"f3c2b172",
   299 => x"4abf97f1",
   300 => x"c29dcf4d",
   301 => x"bf97f2f3",
   302 => x"ca9ac34a",
   303 => x"f3f3c232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97f4f3",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"d2fcc286",
   323 => x"c278c048",
   324 => x"c01ecaf4",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfd0f8c0",
   331 => x"c0f5c249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f8c07ec0",
   336 => x"c249bfcc",
   337 => x"714adcf5",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"d0fbc287",
   343 => x"fcc24dbf",
   344 => x"7ebf9fc8",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bfd0fbc2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"caf4c287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f8c087dc",
   358 => x"c249bfcc",
   359 => x"714adcf5",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"fcc287c8",
   363 => x"78c148d2",
   364 => x"f8c087da",
   365 => x"c249bfd0",
   366 => x"714ac0f5",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97c8fcc2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"c9fcc287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97caf4",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97d5f4",
   387 => x"c0059949",
   388 => x"f4c287cc",
   389 => x"49bf97d6",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97d7f4",
   394 => x"cefcc248",
   395 => x"484c7058",
   396 => x"fcc288c1",
   397 => x"f4c258d2",
   398 => x"49bf97d8",
   399 => x"f4c28175",
   400 => x"4abf97d9",
   401 => x"a17232c8",
   402 => x"dfc0c37e",
   403 => x"c2786e48",
   404 => x"bf97daf4",
   405 => x"58a6c848",
   406 => x"bfd2fcc2",
   407 => x"87d4c202",
   408 => x"bfccf8c0",
   409 => x"dcf5c249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"fcc287f8",
   415 => x"c34cbfca",
   416 => x"c25cf3c0",
   417 => x"bf97eff4",
   418 => x"c231c849",
   419 => x"bf97eef4",
   420 => x"c249a14a",
   421 => x"bf97f0f4",
   422 => x"7232d04a",
   423 => x"f4c249a1",
   424 => x"4abf97f1",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfdfc0c3",
   428 => x"e7c0c381",
   429 => x"f7f4c259",
   430 => x"c84abf97",
   431 => x"f6f4c232",
   432 => x"a24bbf97",
   433 => x"f8f4c24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97f9f4c2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"ebc0c34a",
   440 => x"e7c0c35a",
   441 => x"8ac24abf",
   442 => x"c0c39274",
   443 => x"a17248eb",
   444 => x"87cac178",
   445 => x"97dcf4c2",
   446 => x"31c849bf",
   447 => x"97dbf4c2",
   448 => x"49a14abf",
   449 => x"59dafcc2",
   450 => x"bfd6fcc2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59f3c0c3",
   454 => x"97e1f4c2",
   455 => x"32c84abf",
   456 => x"97e0f4c2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"efc0c382",
   460 => x"e7c0c35a",
   461 => x"c378c048",
   462 => x"7248e3c0",
   463 => x"c0c378a1",
   464 => x"c0c348f3",
   465 => x"c378bfe7",
   466 => x"c348f7c0",
   467 => x"78bfebc0",
   468 => x"bfd2fcc2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"efc0c387",
   473 => x"30c448bf",
   474 => x"fcc27e70",
   475 => x"786e48d6",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bfd2fcc2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c39cffc3",
   488 => x"83bfdfc0",
   489 => x"bfc8f8c0",
   490 => x"87d902ab",
   491 => x"5bccf8c0",
   492 => x"1ecaf4c2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"d2fcc287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81caf4c2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"f4c291c2",
   505 => x"699f81ca",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"d049c11e",
   511 => x"86c487f2",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754adafc",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"cf4966c4",
   527 => x"86c487f2",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"f80e5d5c",
   533 => x"9b4b7186",
   534 => x"c087c505",
   535 => x"87d4c248",
   536 => x"c04da3c8",
   537 => x"0266d87d",
   538 => x"66d887c7",
   539 => x"c505bf97",
   540 => x"c148c087",
   541 => x"66d887fe",
   542 => x"87f2fd49",
   543 => x"026e7e70",
   544 => x"6e87efc1",
   545 => x"6981dc49",
   546 => x"da496e7d",
   547 => x"4ca3c481",
   548 => x"c27c699f",
   549 => x"02bfd2fc",
   550 => x"496e87d0",
   551 => x"699f81d4",
   552 => x"ffc04a49",
   553 => x"32d09aff",
   554 => x"4ac087c2",
   555 => x"6c484972",
   556 => x"c07c7080",
   557 => x"49a3cc7b",
   558 => x"a3d0796c",
   559 => x"c479c049",
   560 => x"78c048a6",
   561 => x"c44aa3d4",
   562 => x"91c84966",
   563 => x"c049a172",
   564 => x"c4796c41",
   565 => x"80c14866",
   566 => x"c458a6c8",
   567 => x"ff04a8b7",
   568 => x"4a6d87e2",
   569 => x"2ac52ac9",
   570 => x"49a3f4c0",
   571 => x"486e7972",
   572 => x"48c087c2",
   573 => x"fbf98ef8",
   574 => x"5b5e0e87",
   575 => x"710e5d5c",
   576 => x"c8f8c04c",
   577 => x"7478ff48",
   578 => x"cac1029c",
   579 => x"49a4c887",
   580 => x"c2c10269",
   581 => x"4a66d087",
   582 => x"d482496c",
   583 => x"66d05aa6",
   584 => x"fcc2b94d",
   585 => x"ff4abfce",
   586 => x"719972ba",
   587 => x"e4c00299",
   588 => x"4ba4c487",
   589 => x"c3f9496b",
   590 => x"c27b7087",
   591 => x"49bfcafc",
   592 => x"7c71816c",
   593 => x"fcc2b975",
   594 => x"ff4abfce",
   595 => x"719972ba",
   596 => x"dcff0599",
   597 => x"f87c7587",
   598 => x"731e87da",
   599 => x"9b4b711e",
   600 => x"c887c702",
   601 => x"056949a3",
   602 => x"48c087c5",
   603 => x"c387ebc0",
   604 => x"4abfe3c0",
   605 => x"6949a3c4",
   606 => x"c289c249",
   607 => x"91bfcafc",
   608 => x"c24aa271",
   609 => x"49bfcefc",
   610 => x"a271996b",
   611 => x"1e66c84a",
   612 => x"e1e94972",
   613 => x"7086c487",
   614 => x"dbf74849",
   615 => x"1e731e87",
   616 => x"029b4b71",
   617 => x"a3c887c7",
   618 => x"c5056949",
   619 => x"c048c087",
   620 => x"c0c387eb",
   621 => x"c44abfe3",
   622 => x"496949a3",
   623 => x"fcc289c2",
   624 => x"7191bfca",
   625 => x"fcc24aa2",
   626 => x"6b49bfce",
   627 => x"4aa27199",
   628 => x"721e66c8",
   629 => x"87d4e549",
   630 => x"497086c4",
   631 => x"87d8f648",
   632 => x"5c5b5e0e",
   633 => x"86f80e5d",
   634 => x"a6c44b71",
   635 => x"c878ff48",
   636 => x"4d6949a3",
   637 => x"a3d44cc0",
   638 => x"c849744a",
   639 => x"49a17291",
   640 => x"66d84969",
   641 => x"70887148",
   642 => x"a966d87e",
   643 => x"6e87ca01",
   644 => x"87c506ad",
   645 => x"6e5ca6c8",
   646 => x"c484c14d",
   647 => x"ff04acb7",
   648 => x"486687d4",
   649 => x"cbf58ef8",
   650 => x"5b5e0e87",
   651 => x"ec0e5d5c",
   652 => x"59a6c886",
   653 => x"c148a6c8",
   654 => x"ffffffff",
   655 => x"80c478ff",
   656 => x"4dc078ff",
   657 => x"66c44cc0",
   658 => x"7483d44b",
   659 => x"7391c849",
   660 => x"4a7549a1",
   661 => x"a27392c8",
   662 => x"6e49697e",
   663 => x"a6d489bf",
   664 => x"05ad7459",
   665 => x"a6d087c6",
   666 => x"78bf6e48",
   667 => x"c04866d0",
   668 => x"cf04a8b7",
   669 => x"4966d087",
   670 => x"03a966c8",
   671 => x"a6d087c6",
   672 => x"59a6cc5c",
   673 => x"b7c484c1",
   674 => x"f9fe04ac",
   675 => x"c485c187",
   676 => x"fe04adb7",
   677 => x"66cc87ee",
   678 => x"f38eec48",
   679 => x"5e0e87d6",
   680 => x"0e5d5c5b",
   681 => x"4b7186f0",
   682 => x"4c66e0c0",
   683 => x"9b732cc9",
   684 => x"87e1c302",
   685 => x"6949a3c8",
   686 => x"87d9c302",
   687 => x"c049a3d0",
   688 => x"6b7966e0",
   689 => x"c302ac7e",
   690 => x"fcc287cb",
   691 => x"ff49bfce",
   692 => x"744a71b9",
   693 => x"6e48719a",
   694 => x"58a6cc98",
   695 => x"c44da3c4",
   696 => x"786d48a6",
   697 => x"05aa66c8",
   698 => x"7b7487c5",
   699 => x"7287d1c2",
   700 => x"fb49731e",
   701 => x"86c487ea",
   702 => x"c0487e70",
   703 => x"d004a8b7",
   704 => x"4aa3d487",
   705 => x"91c8496e",
   706 => x"2149a172",
   707 => x"c77d697b",
   708 => x"cc7bc087",
   709 => x"7d6949a3",
   710 => x"731e66c8",
   711 => x"87c0fb49",
   712 => x"7e7086c4",
   713 => x"49a3f4c0",
   714 => x"6948a6cc",
   715 => x"4866c878",
   716 => x"06a866cc",
   717 => x"486e87c9",
   718 => x"04a8b7c0",
   719 => x"6e87e0c0",
   720 => x"a8b7c048",
   721 => x"87ecc004",
   722 => x"6e4aa3d4",
   723 => x"7291c849",
   724 => x"66c849a1",
   725 => x"70886948",
   726 => x"a966cc49",
   727 => x"7387d506",
   728 => x"87c5fb49",
   729 => x"a3d44970",
   730 => x"7291c84a",
   731 => x"66c849a1",
   732 => x"7966c441",
   733 => x"49748c6b",
   734 => x"f549731e",
   735 => x"86c487fb",
   736 => x"4966e0c0",
   737 => x"0299ffc7",
   738 => x"f4c287cb",
   739 => x"49731eca",
   740 => x"c487c7f7",
   741 => x"ef8ef086",
   742 => x"731e87da",
   743 => x"9b4b711e",
   744 => x"87e4c002",
   745 => x"5bf7c0c3",
   746 => x"8ac24a73",
   747 => x"bfcafcc2",
   748 => x"c0c39249",
   749 => x"7248bfe3",
   750 => x"fbc0c380",
   751 => x"c4487158",
   752 => x"dafcc230",
   753 => x"87edc058",
   754 => x"48f3c0c3",
   755 => x"bfe7c0c3",
   756 => x"f7c0c378",
   757 => x"ebc0c348",
   758 => x"fcc278bf",
   759 => x"c902bfd2",
   760 => x"cafcc287",
   761 => x"31c449bf",
   762 => x"c0c387c7",
   763 => x"c449bfef",
   764 => x"dafcc231",
   765 => x"87c0ee59",
   766 => x"5c5b5e0e",
   767 => x"c04a710e",
   768 => x"029a724b",
   769 => x"da87e1c0",
   770 => x"699f49a2",
   771 => x"d2fcc24b",
   772 => x"87cf02bf",
   773 => x"9f49a2d4",
   774 => x"c04c4969",
   775 => x"d09cffff",
   776 => x"c087c234",
   777 => x"b349744c",
   778 => x"edfd4973",
   779 => x"87c6ed87",
   780 => x"5c5b5e0e",
   781 => x"86f40e5d",
   782 => x"7ec04a71",
   783 => x"d8029a72",
   784 => x"c6f4c287",
   785 => x"c278c048",
   786 => x"c348fef3",
   787 => x"78bff7c0",
   788 => x"48c2f4c2",
   789 => x"bff3c0c3",
   790 => x"e7fcc278",
   791 => x"c250c048",
   792 => x"49bfd6fc",
   793 => x"bfc6f4c2",
   794 => x"03aa714a",
   795 => x"7287c0c4",
   796 => x"0599cf49",
   797 => x"c287e1c0",
   798 => x"c21ecaf4",
   799 => x"49bffef3",
   800 => x"48fef3c2",
   801 => x"7178a1c1",
   802 => x"87eaddff",
   803 => x"f8c086c4",
   804 => x"f4c248c4",
   805 => x"87cc78ca",
   806 => x"bfc4f8c0",
   807 => x"80e0c048",
   808 => x"58c8f8c0",
   809 => x"bfc6f4c2",
   810 => x"c280c148",
   811 => x"2758caf4",
   812 => x"00000e04",
   813 => x"4dbf97bf",
   814 => x"e2c2029d",
   815 => x"ade5c387",
   816 => x"87dbc202",
   817 => x"bfc4f8c0",
   818 => x"49a3cb4b",
   819 => x"accf4c11",
   820 => x"87d2c105",
   821 => x"99df4975",
   822 => x"91cd89c1",
   823 => x"81dafcc2",
   824 => x"124aa3c1",
   825 => x"4aa3c351",
   826 => x"a3c55112",
   827 => x"c751124a",
   828 => x"51124aa3",
   829 => x"124aa3c9",
   830 => x"4aa3ce51",
   831 => x"a3d05112",
   832 => x"d251124a",
   833 => x"51124aa3",
   834 => x"124aa3d4",
   835 => x"4aa3d651",
   836 => x"a3d85112",
   837 => x"dc51124a",
   838 => x"51124aa3",
   839 => x"124aa3de",
   840 => x"c07ec151",
   841 => x"497487f9",
   842 => x"c00599c8",
   843 => x"497487ea",
   844 => x"d00599d0",
   845 => x"0266dc87",
   846 => x"7387cac0",
   847 => x"0f66dc49",
   848 => x"d3029870",
   849 => x"c0056e87",
   850 => x"fcc287c6",
   851 => x"50c048da",
   852 => x"bfc4f8c0",
   853 => x"87e7c248",
   854 => x"48e7fcc2",
   855 => x"c27e50c0",
   856 => x"49bfd6fc",
   857 => x"bfc6f4c2",
   858 => x"04aa714a",
   859 => x"c387c0fc",
   860 => x"05bff7c0",
   861 => x"c287c8c0",
   862 => x"02bfd2fc",
   863 => x"c087fec1",
   864 => x"ff48c8f8",
   865 => x"c2f4c278",
   866 => x"efe749bf",
   867 => x"c2497087",
   868 => x"c459c6f4",
   869 => x"f4c248a6",
   870 => x"c278bfc2",
   871 => x"02bfd2fc",
   872 => x"c487d8c0",
   873 => x"ffcf4966",
   874 => x"99f8ffff",
   875 => x"c5c002a9",
   876 => x"c04dc087",
   877 => x"4dc187e1",
   878 => x"c487dcc0",
   879 => x"ffcf4966",
   880 => x"02a999f8",
   881 => x"c887c8c0",
   882 => x"78c048a6",
   883 => x"c887c5c0",
   884 => x"78c148a6",
   885 => x"754d66c8",
   886 => x"e0c0059d",
   887 => x"4966c487",
   888 => x"fcc289c2",
   889 => x"914abfca",
   890 => x"bfe3c0c3",
   891 => x"fef3c24a",
   892 => x"78a17248",
   893 => x"48c6f4c2",
   894 => x"e2f978c0",
   895 => x"f448c087",
   896 => x"87f0e58e",
   897 => x"00000000",
   898 => x"ffffffff",
   899 => x"00000e14",
   900 => x"00000e1d",
   901 => x"33544146",
   902 => x"20202032",
   903 => x"54414600",
   904 => x"20203631",
   905 => x"ff1e0020",
   906 => x"ffc348d4",
   907 => x"26486878",
   908 => x"d4ff1e4f",
   909 => x"78ffc348",
   910 => x"c848d0ff",
   911 => x"d4ff78e1",
   912 => x"c378d448",
   913 => x"ff48fbc0",
   914 => x"2650bfd4",
   915 => x"d0ff1e4f",
   916 => x"78e0c048",
   917 => x"ff1e4f26",
   918 => x"497087cc",
   919 => x"87c60299",
   920 => x"05a9fbc0",
   921 => x"487187f1",
   922 => x"5e0e4f26",
   923 => x"710e5c5b",
   924 => x"fe4cc04b",
   925 => x"497087f0",
   926 => x"f9c00299",
   927 => x"a9ecc087",
   928 => x"87f2c002",
   929 => x"02a9fbc0",
   930 => x"cc87ebc0",
   931 => x"03acb766",
   932 => x"66d087c7",
   933 => x"7187c202",
   934 => x"02997153",
   935 => x"84c187c2",
   936 => x"7087c3fe",
   937 => x"cd029949",
   938 => x"a9ecc087",
   939 => x"c087c702",
   940 => x"ff05a9fb",
   941 => x"66d087d5",
   942 => x"c087c302",
   943 => x"ecc07b97",
   944 => x"87c405a9",
   945 => x"87c54a74",
   946 => x"0ac04a74",
   947 => x"c248728a",
   948 => x"264d2687",
   949 => x"264b264c",
   950 => x"c9fd1e4f",
   951 => x"c0497087",
   952 => x"04a9b7f0",
   953 => x"f9c087ca",
   954 => x"c301a9b7",
   955 => x"89f0c087",
   956 => x"a9b7c1c1",
   957 => x"c187ca04",
   958 => x"01a9b7da",
   959 => x"f7c087c3",
   960 => x"b7e1c189",
   961 => x"87ca04a9",
   962 => x"a9b7fac1",
   963 => x"c087c301",
   964 => x"487189fd",
   965 => x"5e0e4f26",
   966 => x"710e5c5b",
   967 => x"4cd4ff4a",
   968 => x"eac04972",
   969 => x"9b4b7087",
   970 => x"c187c202",
   971 => x"48d0ff8b",
   972 => x"c178c5c8",
   973 => x"49737cd5",
   974 => x"f2c231c6",
   975 => x"4abf97f3",
   976 => x"70b07148",
   977 => x"48d0ff7c",
   978 => x"487378c4",
   979 => x"0e87c4fe",
   980 => x"5d5c5b5e",
   981 => x"7186f80e",
   982 => x"fb7ec04c",
   983 => x"4bc087d3",
   984 => x"97fcffc0",
   985 => x"a9c049bf",
   986 => x"fb87cf04",
   987 => x"83c187e8",
   988 => x"97fcffc0",
   989 => x"06ab49bf",
   990 => x"ffc087f1",
   991 => x"02bf97fc",
   992 => x"e1fa87cf",
   993 => x"99497087",
   994 => x"c087c602",
   995 => x"f105a9ec",
   996 => x"fa4bc087",
   997 => x"4d7087d0",
   998 => x"c887cbfa",
   999 => x"c5fa58a6",
  1000 => x"c14a7087",
  1001 => x"49a4c883",
  1002 => x"ad496997",
  1003 => x"c087c702",
  1004 => x"c005adff",
  1005 => x"a4c987e7",
  1006 => x"49699749",
  1007 => x"02a966c4",
  1008 => x"c04887c7",
  1009 => x"d405a8ff",
  1010 => x"49a4ca87",
  1011 => x"aa496997",
  1012 => x"c087c602",
  1013 => x"c405aaff",
  1014 => x"d07ec187",
  1015 => x"adecc087",
  1016 => x"c087c602",
  1017 => x"c405adfb",
  1018 => x"c14bc087",
  1019 => x"fe026e7e",
  1020 => x"d8f987e1",
  1021 => x"f8487387",
  1022 => x"87d5fb8e",
  1023 => x"5b5e0e00",
  1024 => x"1e0e5d5c",
  1025 => x"4cc04b71",
  1026 => x"c004ab4d",
  1027 => x"fdc087e8",
  1028 => x"9d751ecf",
  1029 => x"c087c402",
  1030 => x"c187c24a",
  1031 => x"f049724a",
  1032 => x"86c487ce",
  1033 => x"84c17e70",
  1034 => x"87c2056e",
  1035 => x"85c14c73",
  1036 => x"ff06ac73",
  1037 => x"486e87d8",
  1038 => x"264d2626",
  1039 => x"264b264c",
  1040 => x"5b5e0e4f",
  1041 => x"1e0e5d5c",
  1042 => x"de494c71",
  1043 => x"d5c1c391",
  1044 => x"9785714d",
  1045 => x"ddc1026d",
  1046 => x"c0c1c387",
  1047 => x"82744abf",
  1048 => x"d8fe4972",
  1049 => x"6e7e7087",
  1050 => x"87f3c002",
  1051 => x"4bc8c1c3",
  1052 => x"49cb4a6e",
  1053 => x"87f0c0ff",
  1054 => x"93cb4b74",
  1055 => x"83f5e3c1",
  1056 => x"c2c183c4",
  1057 => x"49747bfa",
  1058 => x"87ebd4c1",
  1059 => x"c1c37b75",
  1060 => x"49bf97d4",
  1061 => x"c8c1c31e",
  1062 => x"d8efc149",
  1063 => x"7486c487",
  1064 => x"d2d4c149",
  1065 => x"c149c087",
  1066 => x"c387f1d5",
  1067 => x"c048fcc0",
  1068 => x"dd49c178",
  1069 => x"fd2687d0",
  1070 => x"6f4c87ff",
  1071 => x"6e696461",
  1072 => x"2e2e2e67",
  1073 => x"5b5e0e00",
  1074 => x"4b710e5c",
  1075 => x"c0c1c34a",
  1076 => x"497282bf",
  1077 => x"7087e6fc",
  1078 => x"c4029c4c",
  1079 => x"d7ec4987",
  1080 => x"c0c1c387",
  1081 => x"c178c048",
  1082 => x"87dadc49",
  1083 => x"0e87ccfd",
  1084 => x"5d5c5b5e",
  1085 => x"c286f40e",
  1086 => x"c04dcaf4",
  1087 => x"48a6c44c",
  1088 => x"c1c378c0",
  1089 => x"c049bfc0",
  1090 => x"c1c106a9",
  1091 => x"caf4c287",
  1092 => x"c0029848",
  1093 => x"fdc087f8",
  1094 => x"66c81ecf",
  1095 => x"c487c702",
  1096 => x"78c048a6",
  1097 => x"a6c487c5",
  1098 => x"c478c148",
  1099 => x"ffeb4966",
  1100 => x"7086c487",
  1101 => x"c484c14d",
  1102 => x"80c14866",
  1103 => x"c358a6c8",
  1104 => x"49bfc0c1",
  1105 => x"87c603ac",
  1106 => x"ff059d75",
  1107 => x"4cc087c8",
  1108 => x"c3029d75",
  1109 => x"fdc087e0",
  1110 => x"66c81ecf",
  1111 => x"cc87c702",
  1112 => x"78c048a6",
  1113 => x"a6cc87c5",
  1114 => x"cc78c148",
  1115 => x"ffea4966",
  1116 => x"7086c487",
  1117 => x"c2026e7e",
  1118 => x"496e87e9",
  1119 => x"699781cb",
  1120 => x"0299d049",
  1121 => x"c187d6c1",
  1122 => x"744ac5c3",
  1123 => x"c191cb49",
  1124 => x"7281f5e3",
  1125 => x"c381c879",
  1126 => x"497451ff",
  1127 => x"c1c391de",
  1128 => x"85714dd5",
  1129 => x"7d97c1c2",
  1130 => x"c049a5c1",
  1131 => x"fcc251e0",
  1132 => x"02bf97da",
  1133 => x"84c187d2",
  1134 => x"c24ba5c2",
  1135 => x"db4adafc",
  1136 => x"e3fbfe49",
  1137 => x"87dbc187",
  1138 => x"c049a5cd",
  1139 => x"c284c151",
  1140 => x"4a6e4ba5",
  1141 => x"fbfe49cb",
  1142 => x"c6c187ce",
  1143 => x"c1c1c187",
  1144 => x"cb49744a",
  1145 => x"f5e3c191",
  1146 => x"c2797281",
  1147 => x"bf97dafc",
  1148 => x"7487d802",
  1149 => x"c191de49",
  1150 => x"d5c1c384",
  1151 => x"c283714b",
  1152 => x"dd4adafc",
  1153 => x"dffafe49",
  1154 => x"7487d887",
  1155 => x"c393de4b",
  1156 => x"cb83d5c1",
  1157 => x"51c049a3",
  1158 => x"6e7384c1",
  1159 => x"fe49cb4a",
  1160 => x"c487c5fa",
  1161 => x"80c14866",
  1162 => x"c758a6c8",
  1163 => x"c5c003ac",
  1164 => x"fc056e87",
  1165 => x"487487e0",
  1166 => x"fcf78ef4",
  1167 => x"1e731e87",
  1168 => x"cb494b71",
  1169 => x"f5e3c191",
  1170 => x"4aa1c881",
  1171 => x"48f3f2c2",
  1172 => x"a1c95012",
  1173 => x"fcffc04a",
  1174 => x"ca501248",
  1175 => x"d4c1c381",
  1176 => x"c3501148",
  1177 => x"bf97d4c1",
  1178 => x"49c01e49",
  1179 => x"87c5e8c1",
  1180 => x"48fcc0c3",
  1181 => x"49c178de",
  1182 => x"2687cbd6",
  1183 => x"1e87fef6",
  1184 => x"cb494a71",
  1185 => x"f5e3c191",
  1186 => x"1181c881",
  1187 => x"c0c1c348",
  1188 => x"c0c1c358",
  1189 => x"c178c048",
  1190 => x"87ead549",
  1191 => x"c01e4f26",
  1192 => x"f7cdc149",
  1193 => x"1e4f2687",
  1194 => x"d2029971",
  1195 => x"cae5c187",
  1196 => x"f750c048",
  1197 => x"ffc9c180",
  1198 => x"eee3c140",
  1199 => x"c187ce78",
  1200 => x"c148c6e5",
  1201 => x"fc78e7e3",
  1202 => x"decac180",
  1203 => x"0e4f2678",
  1204 => x"0e5c5b5e",
  1205 => x"cb4a4c71",
  1206 => x"f5e3c192",
  1207 => x"49a2c882",
  1208 => x"974ba2c9",
  1209 => x"971e4b6b",
  1210 => x"ca1e4969",
  1211 => x"c0491282",
  1212 => x"c087f0f6",
  1213 => x"87ced449",
  1214 => x"cac14974",
  1215 => x"8ef887f9",
  1216 => x"1e87f8f4",
  1217 => x"4b711e73",
  1218 => x"87c3ff49",
  1219 => x"fefe4973",
  1220 => x"c149c087",
  1221 => x"f487c5cc",
  1222 => x"731e87e3",
  1223 => x"c64b711e",
  1224 => x"db024aa3",
  1225 => x"028ac187",
  1226 => x"028a87d6",
  1227 => x"8a87dac1",
  1228 => x"87fcc002",
  1229 => x"e1c0028a",
  1230 => x"cb028a87",
  1231 => x"87dbc187",
  1232 => x"fafc49c7",
  1233 => x"87dec187",
  1234 => x"bfc0c1c3",
  1235 => x"87cbc102",
  1236 => x"c388c148",
  1237 => x"c158c4c1",
  1238 => x"c1c387c1",
  1239 => x"c002bfc4",
  1240 => x"c1c387f9",
  1241 => x"c148bfc0",
  1242 => x"c4c1c380",
  1243 => x"87ebc058",
  1244 => x"bfc0c1c3",
  1245 => x"c389c649",
  1246 => x"c059c4c1",
  1247 => x"da03a9b7",
  1248 => x"c0c1c387",
  1249 => x"d278c048",
  1250 => x"c4c1c387",
  1251 => x"87cb02bf",
  1252 => x"bfc0c1c3",
  1253 => x"c380c648",
  1254 => x"c058c4c1",
  1255 => x"87e6d149",
  1256 => x"c8c14973",
  1257 => x"d4f287d1",
  1258 => x"5b5e0e87",
  1259 => x"4c710e5c",
  1260 => x"741e66cc",
  1261 => x"c193cb4b",
  1262 => x"c483f5e3",
  1263 => x"496a4aa3",
  1264 => x"87f4f3fe",
  1265 => x"7bfdc8c1",
  1266 => x"d449a3c8",
  1267 => x"a3c95166",
  1268 => x"5166d849",
  1269 => x"dc49a3ca",
  1270 => x"f1265166",
  1271 => x"5e0e87dd",
  1272 => x"0e5d5c5b",
  1273 => x"d886d0ff",
  1274 => x"a6c459a6",
  1275 => x"c478c048",
  1276 => x"66c4c180",
  1277 => x"c180c478",
  1278 => x"c180c478",
  1279 => x"c4c1c378",
  1280 => x"c378c148",
  1281 => x"48bffcc0",
  1282 => x"cb05a8de",
  1283 => x"87dff387",
  1284 => x"a6c84970",
  1285 => x"87f7ce59",
  1286 => x"e887d6e8",
  1287 => x"c5e887f8",
  1288 => x"c04c7087",
  1289 => x"c102acfb",
  1290 => x"66d487d0",
  1291 => x"87c2c105",
  1292 => x"c11e1ec0",
  1293 => x"e8e5c11e",
  1294 => x"fd49c01e",
  1295 => x"d0c187eb",
  1296 => x"82c44a66",
  1297 => x"81c7496a",
  1298 => x"1ec15174",
  1299 => x"496a1ed8",
  1300 => x"d5e881c8",
  1301 => x"c186d887",
  1302 => x"c04866c4",
  1303 => x"87c701a8",
  1304 => x"c148a6c4",
  1305 => x"c187ce78",
  1306 => x"c14866c4",
  1307 => x"58a6cc88",
  1308 => x"e1e787c3",
  1309 => x"48a6cc87",
  1310 => x"9c7478c2",
  1311 => x"87cbcd02",
  1312 => x"c14866c4",
  1313 => x"03a866c8",
  1314 => x"d887c0cd",
  1315 => x"78c048a6",
  1316 => x"7087d3e6",
  1317 => x"acd0c14c",
  1318 => x"87d6c205",
  1319 => x"e87e66d8",
  1320 => x"497087f7",
  1321 => x"e559a6dc",
  1322 => x"4c7087fc",
  1323 => x"05acecc0",
  1324 => x"c487eac1",
  1325 => x"91cb4966",
  1326 => x"8166c0c1",
  1327 => x"6a4aa1c4",
  1328 => x"4aa1c84d",
  1329 => x"c15266d8",
  1330 => x"e579ffc9",
  1331 => x"4c7087d8",
  1332 => x"87d8029c",
  1333 => x"02acfbc0",
  1334 => x"557487d2",
  1335 => x"7087c7e5",
  1336 => x"c7029c4c",
  1337 => x"acfbc087",
  1338 => x"87eeff05",
  1339 => x"c255e0c0",
  1340 => x"97c055c1",
  1341 => x"4966d47d",
  1342 => x"db05a96e",
  1343 => x"4866c487",
  1344 => x"04a866c8",
  1345 => x"66c487ca",
  1346 => x"c880c148",
  1347 => x"87c858a6",
  1348 => x"c14866c8",
  1349 => x"58a6cc88",
  1350 => x"7087cbe4",
  1351 => x"acd0c14c",
  1352 => x"d087c805",
  1353 => x"80c14866",
  1354 => x"c158a6d4",
  1355 => x"fd02acd0",
  1356 => x"a6dc87ea",
  1357 => x"7866d448",
  1358 => x"dc4866d8",
  1359 => x"c905a866",
  1360 => x"e0c087db",
  1361 => x"f0c048a6",
  1362 => x"cc80c478",
  1363 => x"80c47866",
  1364 => x"747e78c0",
  1365 => x"88fbc048",
  1366 => x"58a6f0c0",
  1367 => x"c8029870",
  1368 => x"cb4887d6",
  1369 => x"a6f0c088",
  1370 => x"02987058",
  1371 => x"4887e9c0",
  1372 => x"f0c088c9",
  1373 => x"987058a6",
  1374 => x"87e1c302",
  1375 => x"c088c448",
  1376 => x"7058a6f0",
  1377 => x"87de0298",
  1378 => x"c088c148",
  1379 => x"7058a6f0",
  1380 => x"c8c30298",
  1381 => x"87dac787",
  1382 => x"48a6e0c0",
  1383 => x"66cc78c0",
  1384 => x"d080c148",
  1385 => x"fde158a6",
  1386 => x"c04c7087",
  1387 => x"d502acec",
  1388 => x"66e0c087",
  1389 => x"c087c602",
  1390 => x"c95ca6e4",
  1391 => x"c0487487",
  1392 => x"e8c088f0",
  1393 => x"ecc058a6",
  1394 => x"87cc02ac",
  1395 => x"7087d7e1",
  1396 => x"acecc04c",
  1397 => x"87f4ff05",
  1398 => x"1e66e0c0",
  1399 => x"1e4966d4",
  1400 => x"1e66ecc0",
  1401 => x"1ee8e5c1",
  1402 => x"f64966d4",
  1403 => x"1ec087fb",
  1404 => x"66dc1eca",
  1405 => x"c191cb49",
  1406 => x"d88166d8",
  1407 => x"a1c448a6",
  1408 => x"bf66d878",
  1409 => x"87e2e149",
  1410 => x"b7c086d8",
  1411 => x"c7c106a8",
  1412 => x"de1ec187",
  1413 => x"bf66c81e",
  1414 => x"87cee149",
  1415 => x"497086c8",
  1416 => x"8808c048",
  1417 => x"58a6e4c0",
  1418 => x"06a8b7c0",
  1419 => x"c087e9c0",
  1420 => x"dd4866e0",
  1421 => x"df03a8b7",
  1422 => x"49bf6e87",
  1423 => x"8166e0c0",
  1424 => x"6651e0c0",
  1425 => x"6e81c149",
  1426 => x"c1c281bf",
  1427 => x"66e0c051",
  1428 => x"6e81c249",
  1429 => x"51c081bf",
  1430 => x"dbc47ec1",
  1431 => x"87f9e187",
  1432 => x"58a6e4c0",
  1433 => x"c087f2e1",
  1434 => x"c058a6e8",
  1435 => x"c005a8ec",
  1436 => x"e4c087cb",
  1437 => x"e0c048a6",
  1438 => x"c4c07866",
  1439 => x"e5deff87",
  1440 => x"4966c487",
  1441 => x"c0c191cb",
  1442 => x"80714866",
  1443 => x"496e7e70",
  1444 => x"4a6e81c8",
  1445 => x"e0c082ca",
  1446 => x"e4c05266",
  1447 => x"82c14a66",
  1448 => x"8a66e0c0",
  1449 => x"307248c1",
  1450 => x"8ac14a70",
  1451 => x"97799772",
  1452 => x"c01e4969",
  1453 => x"c04966e4",
  1454 => x"c487eae6",
  1455 => x"a6f0c086",
  1456 => x"c4496e58",
  1457 => x"dc4d6981",
  1458 => x"66d84866",
  1459 => x"c8c002a8",
  1460 => x"48a6d887",
  1461 => x"c5c078c0",
  1462 => x"48a6d887",
  1463 => x"66d878c1",
  1464 => x"1ee0c01e",
  1465 => x"deff4975",
  1466 => x"86c887c0",
  1467 => x"b7c04c70",
  1468 => x"d4c106ac",
  1469 => x"c0857487",
  1470 => x"897449e0",
  1471 => x"e0c14b75",
  1472 => x"fe714ac3",
  1473 => x"c287e1e6",
  1474 => x"66e8c085",
  1475 => x"c080c148",
  1476 => x"c058a6ec",
  1477 => x"c14966ec",
  1478 => x"02a97081",
  1479 => x"d887c8c0",
  1480 => x"78c048a6",
  1481 => x"d887c5c0",
  1482 => x"78c148a6",
  1483 => x"c21e66d8",
  1484 => x"e0c049a4",
  1485 => x"70887148",
  1486 => x"49751e49",
  1487 => x"87eadcff",
  1488 => x"b7c086c8",
  1489 => x"c0ff01a8",
  1490 => x"66e8c087",
  1491 => x"87d1c002",
  1492 => x"81c9496e",
  1493 => x"5166e8c0",
  1494 => x"cbc1486e",
  1495 => x"ccc078cf",
  1496 => x"c9496e87",
  1497 => x"6e51c281",
  1498 => x"c3ccc148",
  1499 => x"c07ec178",
  1500 => x"dbff87c6",
  1501 => x"4c7087e0",
  1502 => x"f5c0026e",
  1503 => x"4866c487",
  1504 => x"04a866c8",
  1505 => x"c487cbc0",
  1506 => x"80c14866",
  1507 => x"c058a6c8",
  1508 => x"66c887e0",
  1509 => x"cc88c148",
  1510 => x"d5c058a6",
  1511 => x"acc6c187",
  1512 => x"87c8c005",
  1513 => x"c14866cc",
  1514 => x"58a6d080",
  1515 => x"87e6daff",
  1516 => x"66d04c70",
  1517 => x"d480c148",
  1518 => x"9c7458a6",
  1519 => x"87cbc002",
  1520 => x"c14866c4",
  1521 => x"04a866c8",
  1522 => x"ff87c0f3",
  1523 => x"c487fed9",
  1524 => x"a8c74866",
  1525 => x"87e5c003",
  1526 => x"48c4c1c3",
  1527 => x"66c478c0",
  1528 => x"c191cb49",
  1529 => x"c48166c0",
  1530 => x"4a6a4aa1",
  1531 => x"c47952c0",
  1532 => x"80c14866",
  1533 => x"c758a6c8",
  1534 => x"dbff04a8",
  1535 => x"8ed0ff87",
  1536 => x"3a87f6e0",
  1537 => x"731e0020",
  1538 => x"9b4b711e",
  1539 => x"c387c602",
  1540 => x"c048c0c1",
  1541 => x"c31ec778",
  1542 => x"49bfc0c1",
  1543 => x"f5e3c11e",
  1544 => x"fcc0c31e",
  1545 => x"f5ee49bf",
  1546 => x"c386cc87",
  1547 => x"49bffcc0",
  1548 => x"7387f4e9",
  1549 => x"87c8029b",
  1550 => x"49f5e3c1",
  1551 => x"87c9f7c0",
  1552 => x"87f9dfff",
  1553 => x"f3f2c21e",
  1554 => x"c150c048",
  1555 => x"49bfd8e5",
  1556 => x"87f4ccc1",
  1557 => x"4f2648c0",
  1558 => x"87dfcd1e",
  1559 => x"e5fe49c1",
  1560 => x"d6e9fe87",
  1561 => x"02987087",
  1562 => x"f2fe87cd",
  1563 => x"987087d3",
  1564 => x"c187c402",
  1565 => x"c087c24a",
  1566 => x"059a724a",
  1567 => x"1ec087ce",
  1568 => x"49e8e2c1",
  1569 => x"87dec2c1",
  1570 => x"87fe86c4",
  1571 => x"e2c11ec0",
  1572 => x"c2c149f3",
  1573 => x"1ec087d0",
  1574 => x"7087e9fe",
  1575 => x"c5c2c149",
  1576 => x"87e2c387",
  1577 => x"4f268ef8",
  1578 => x"66204453",
  1579 => x"656c6961",
  1580 => x"42002e64",
  1581 => x"69746f6f",
  1582 => x"2e2e676e",
  1583 => x"c01e002e",
  1584 => x"87ced549",
  1585 => x"87e1f9c0",
  1586 => x"87d0c5c1",
  1587 => x"4f2687f1",
  1588 => x"c0c1c31e",
  1589 => x"c378c048",
  1590 => x"c048fcc0",
  1591 => x"87f8fd78",
  1592 => x"c087dbff",
  1593 => x"804f2648",
  1594 => x"69784520",
  1595 => x"20800074",
  1596 => x"6b636142",
  1597 => x"00127f00",
  1598 => x"00305500",
  1599 => x"00000000",
  1600 => x"0000127f",
  1601 => x"00003073",
  1602 => x"7f000000",
  1603 => x"91000012",
  1604 => x"00000030",
  1605 => x"127f0000",
  1606 => x"30af0000",
  1607 => x"00000000",
  1608 => x"00127f00",
  1609 => x"0030cd00",
  1610 => x"00000000",
  1611 => x"0000127f",
  1612 => x"000030eb",
  1613 => x"7f000000",
  1614 => x"09000012",
  1615 => x"00000031",
  1616 => x"127f0000",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"00131a00",
  1620 => x"00000000",
  1621 => x"00000000",
  1622 => x"0000195c",
  1623 => x"544f4f42",
  1624 => x"20202020",
  1625 => x"004d4f52",
  1626 => x"64616f4c",
  1627 => x"002e2a20",
  1628 => x"48f0fe1e",
  1629 => x"09cd78c0",
  1630 => x"4f260979",
  1631 => x"f0fe1e1e",
  1632 => x"26487ebf",
  1633 => x"fe1e4f26",
  1634 => x"78c148f0",
  1635 => x"fe1e4f26",
  1636 => x"78c048f0",
  1637 => x"711e4f26",
  1638 => x"7a97c04a",
  1639 => x"c049a2c1",
  1640 => x"49a2ca51",
  1641 => x"a2cb51c0",
  1642 => x"2651c049",
  1643 => x"5b5e0e4f",
  1644 => x"86f00e5c",
  1645 => x"a4ca4c71",
  1646 => x"7e699749",
  1647 => x"974ba4cb",
  1648 => x"a6c8486b",
  1649 => x"cc80c158",
  1650 => x"98c758a6",
  1651 => x"6e58a6d0",
  1652 => x"a866cc48",
  1653 => x"9787db05",
  1654 => x"6b977e69",
  1655 => x"58a6c848",
  1656 => x"a6cc80c1",
  1657 => x"d098c758",
  1658 => x"486e58a6",
  1659 => x"02a866cc",
  1660 => x"d9fe87e5",
  1661 => x"4aa4cc87",
  1662 => x"72496b97",
  1663 => x"66dc49a1",
  1664 => x"7e6b9751",
  1665 => x"80c1486e",
  1666 => x"c758a6c8",
  1667 => x"58a6cc98",
  1668 => x"c37b9770",
  1669 => x"edfd87d2",
  1670 => x"c28ef087",
  1671 => x"264d2687",
  1672 => x"264b264c",
  1673 => x"5b5e0e4f",
  1674 => x"f40e5d5c",
  1675 => x"974d7186",
  1676 => x"a5c17e6d",
  1677 => x"486c974c",
  1678 => x"6e58a6c8",
  1679 => x"a866c448",
  1680 => x"ff87c505",
  1681 => x"87e6c048",
  1682 => x"c287c3fd",
  1683 => x"6c9749a5",
  1684 => x"4ba3714b",
  1685 => x"974b6b97",
  1686 => x"486e7e6c",
  1687 => x"a6c880c1",
  1688 => x"cc98c758",
  1689 => x"977058a6",
  1690 => x"87dafc7c",
  1691 => x"8ef44873",
  1692 => x"0e87eafe",
  1693 => x"0e5c5b5e",
  1694 => x"4c7186f4",
  1695 => x"c34a66d8",
  1696 => x"a4c29aff",
  1697 => x"496c974b",
  1698 => x"7249a173",
  1699 => x"7e6c9751",
  1700 => x"80c1486e",
  1701 => x"c758a6c8",
  1702 => x"58a6cc98",
  1703 => x"8ef45470",
  1704 => x"1e87fcfd",
  1705 => x"699786f0",
  1706 => x"4aa1c17e",
  1707 => x"c8486a97",
  1708 => x"486e58a6",
  1709 => x"a8b766c4",
  1710 => x"9787d304",
  1711 => x"6a977e69",
  1712 => x"58a6c848",
  1713 => x"66c4486e",
  1714 => x"58a6cc88",
  1715 => x"7e1187d6",
  1716 => x"80c8486e",
  1717 => x"481258a6",
  1718 => x"c458a6cc",
  1719 => x"66c84866",
  1720 => x"58a6d088",
  1721 => x"4f268ef0",
  1722 => x"f41e731e",
  1723 => x"87defa86",
  1724 => x"494bbfe0",
  1725 => x"99c0e0c0",
  1726 => x"7387cb02",
  1727 => x"e7c4c31e",
  1728 => x"87effd49",
  1729 => x"497386c4",
  1730 => x"0299c0d0",
  1731 => x"c387c0c1",
  1732 => x"bf97f1c4",
  1733 => x"f2c4c37e",
  1734 => x"c848bf97",
  1735 => x"486e58a6",
  1736 => x"02a866c4",
  1737 => x"c387e8c0",
  1738 => x"bf97f1c4",
  1739 => x"f3c4c349",
  1740 => x"e0481181",
  1741 => x"c4c37808",
  1742 => x"7ebf97f1",
  1743 => x"80c1486e",
  1744 => x"c758a6c8",
  1745 => x"58a6cc98",
  1746 => x"48f1c4c3",
  1747 => x"e45066c8",
  1748 => x"c0494bbf",
  1749 => x"0299c0e0",
  1750 => x"1e7387cb",
  1751 => x"49fbc4c3",
  1752 => x"c487d0fc",
  1753 => x"d0497386",
  1754 => x"c10299c0",
  1755 => x"c5c387c0",
  1756 => x"7ebf97c5",
  1757 => x"97c6c5c3",
  1758 => x"a6c848bf",
  1759 => x"c4486e58",
  1760 => x"c002a866",
  1761 => x"c5c387e8",
  1762 => x"49bf97c5",
  1763 => x"81c7c5c3",
  1764 => x"08e44811",
  1765 => x"c5c5c378",
  1766 => x"6e7ebf97",
  1767 => x"c880c148",
  1768 => x"98c758a6",
  1769 => x"c358a6cc",
  1770 => x"c848c5c5",
  1771 => x"cbf75066",
  1772 => x"f77e7087",
  1773 => x"8ef487d0",
  1774 => x"1e87e6f9",
  1775 => x"49e7c4c3",
  1776 => x"c387d3f7",
  1777 => x"f749fbc4",
  1778 => x"ebc187cc",
  1779 => x"dff649e8",
  1780 => x"87d9c587",
  1781 => x"5e0e4f26",
  1782 => x"0e5d5c5b",
  1783 => x"bfecc5c3",
  1784 => x"eaf0c14a",
  1785 => x"724c49bf",
  1786 => x"f64d71bc",
  1787 => x"4bc087e0",
  1788 => x"99d04974",
  1789 => x"7587d502",
  1790 => x"7199d049",
  1791 => x"c11ec01e",
  1792 => x"734afcf6",
  1793 => x"c0491282",
  1794 => x"86c887e4",
  1795 => x"832d2cc1",
  1796 => x"ff04abc8",
  1797 => x"edf587da",
  1798 => x"eaf0c187",
  1799 => x"ecc5c348",
  1800 => x"4d2678bf",
  1801 => x"4b264c26",
  1802 => x"00004f26",
  1803 => x"ff1e0000",
  1804 => x"e1c848d0",
  1805 => x"48d4ff78",
  1806 => x"66c478c5",
  1807 => x"c387c302",
  1808 => x"66c878e0",
  1809 => x"ff87c602",
  1810 => x"f0c348d4",
  1811 => x"48d4ff78",
  1812 => x"d0ff7871",
  1813 => x"78e1c848",
  1814 => x"2678e0c0",
  1815 => x"5b5e0e4f",
  1816 => x"4c710e5c",
  1817 => x"49e7c4c3",
  1818 => x"7087faf6",
  1819 => x"aab7c04a",
  1820 => x"87e3c204",
  1821 => x"05aae0c3",
  1822 => x"f4c187c9",
  1823 => x"78c148e0",
  1824 => x"c387d4c2",
  1825 => x"c905aaf0",
  1826 => x"dcf4c187",
  1827 => x"c178c148",
  1828 => x"f4c187f5",
  1829 => x"c702bfe0",
  1830 => x"c24b7287",
  1831 => x"87c2b3c0",
  1832 => x"9c744b72",
  1833 => x"c187d105",
  1834 => x"1ebfdcf4",
  1835 => x"bfe0f4c1",
  1836 => x"fd49721e",
  1837 => x"86c887f8",
  1838 => x"bfdcf4c1",
  1839 => x"87e0c002",
  1840 => x"b7c44973",
  1841 => x"f5c19129",
  1842 => x"4a7381fc",
  1843 => x"92c29acf",
  1844 => x"307248c1",
  1845 => x"baff4a70",
  1846 => x"98694872",
  1847 => x"87db7970",
  1848 => x"b7c44973",
  1849 => x"f5c19129",
  1850 => x"4a7381fc",
  1851 => x"92c29acf",
  1852 => x"307248c3",
  1853 => x"69484a70",
  1854 => x"c17970b0",
  1855 => x"c048e0f4",
  1856 => x"dcf4c178",
  1857 => x"c378c048",
  1858 => x"f449e7c4",
  1859 => x"4a7087d7",
  1860 => x"03aab7c0",
  1861 => x"c087ddfd",
  1862 => x"87c8fc48",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"494a711e",
  1866 => x"2687f2fc",
  1867 => x"4ac01e4f",
  1868 => x"91c44972",
  1869 => x"81fcf5c1",
  1870 => x"82c179c0",
  1871 => x"04aab7d0",
  1872 => x"4f2687ee",
  1873 => x"5c5b5e0e",
  1874 => x"4d710e5d",
  1875 => x"7587fff0",
  1876 => x"2ab7c44a",
  1877 => x"fcf5c192",
  1878 => x"cf4c7582",
  1879 => x"6a94c29c",
  1880 => x"2b744b49",
  1881 => x"48c29bc3",
  1882 => x"4c703074",
  1883 => x"4874bcff",
  1884 => x"7a709871",
  1885 => x"7387cff0",
  1886 => x"87e6fa48",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"25261e16",
  1904 => x"3e3d362e",
  1905 => x"711e731e",
  1906 => x"fbc4c34b",
  1907 => x"87d5f149",
  1908 => x"c41e4970",
  1909 => x"87c4c849",
  1910 => x"c4c386c4",
  1911 => x"c4f149fb",
  1912 => x"ff497087",
  1913 => x"787148d4",
  1914 => x"49fbc4c3",
  1915 => x"7087f6f0",
  1916 => x"48d4ff49",
  1917 => x"d0ff7871",
  1918 => x"78e0c048",
  1919 => x"c705abc4",
  1920 => x"fbc4c387",
  1921 => x"87ddf049",
  1922 => x"4d2687c4",
  1923 => x"4b264c26",
  1924 => x"5e0e4f26",
  1925 => x"0e5d5c5b",
  1926 => x"029a4a71",
  1927 => x"fec187c6",
  1928 => x"78c048ed",
  1929 => x"bfedfec1",
  1930 => x"87c6c105",
  1931 => x"49fbc4c3",
  1932 => x"c087f2ef",
  1933 => x"cd04a8b7",
  1934 => x"fbc4c387",
  1935 => x"87e5ef49",
  1936 => x"03a8b7c0",
  1937 => x"fec187f3",
  1938 => x"c149bfed",
  1939 => x"c148edfe",
  1940 => x"fec178a1",
  1941 => x"481181fd",
  1942 => x"58f5fec1",
  1943 => x"48f5fec1",
  1944 => x"f2c078c0",
  1945 => x"daecc049",
  1946 => x"c3497087",
  1947 => x"c459d3c5",
  1948 => x"fec187f8",
  1949 => x"c102bff5",
  1950 => x"c4c387f2",
  1951 => x"e4ee49fb",
  1952 => x"a8b7c087",
  1953 => x"c187cd04",
  1954 => x"48bff5fe",
  1955 => x"fec188c1",
  1956 => x"87db58f9",
  1957 => x"bfcfc5c3",
  1958 => x"f2ebc049",
  1959 => x"02987087",
  1960 => x"c4c387cd",
  1961 => x"edeb49fb",
  1962 => x"edfec187",
  1963 => x"c178c048",
  1964 => x"05bff1fe",
  1965 => x"c187f3c3",
  1966 => x"05bff5fe",
  1967 => x"c187ebc3",
  1968 => x"49bfedfe",
  1969 => x"48edfec1",
  1970 => x"c178a1c1",
  1971 => x"1181fdfe",
  1972 => x"c0c2494b",
  1973 => x"ccc00299",
  1974 => x"c1487387",
  1975 => x"fec198ff",
  1976 => x"c5c358f9",
  1977 => x"f5fec187",
  1978 => x"87fec25b",
  1979 => x"bff1fec1",
  1980 => x"87dbc102",
  1981 => x"bfcfc5c3",
  1982 => x"d2eac049",
  1983 => x"02987087",
  1984 => x"c187e7c2",
  1985 => x"49bfedfe",
  1986 => x"48edfec1",
  1987 => x"c178a1c1",
  1988 => x"9781fdfe",
  1989 => x"c31e4969",
  1990 => x"ea49fbc4",
  1991 => x"86c487cf",
  1992 => x"bff1fec1",
  1993 => x"c189c149",
  1994 => x"c159f5fe",
  1995 => x"c148f5fe",
  1996 => x"02997178",
  1997 => x"c087c6c0",
  1998 => x"c3c04cf2",
  1999 => x"4cdcd787",
  2000 => x"e8c04974",
  2001 => x"497087fd",
  2002 => x"59d3c5c3",
  2003 => x"c387dbc1",
  2004 => x"ed49fbc4",
  2005 => x"4b7087cd",
  2006 => x"eec0029b",
  2007 => x"f9fec187",
  2008 => x"03abb7bf",
  2009 => x"c387e4c0",
  2010 => x"49bfcfc5",
  2011 => x"87dfe8c0",
  2012 => x"c0029870",
  2013 => x"48c787f4",
  2014 => x"bff9fec1",
  2015 => x"fdfec188",
  2016 => x"fbc4c358",
  2017 => x"87cee849",
  2018 => x"d787dfc0",
  2019 => x"e7c049dc",
  2020 => x"497087f1",
  2021 => x"59d3c5c3",
  2022 => x"bff9fec1",
  2023 => x"04abb74a",
  2024 => x"4987c7c0",
  2025 => x"fe87ddf8",
  2026 => x"ddf987e5",
  2027 => x"00000087",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000400",
  2031 => x"82ff0100",
  2032 => x"f3c8f308",
  2033 => x"f250f364",
  2034 => x"f4018101",
  2035 => x"d0ff1e00",
  2036 => x"78e1c848",
  2037 => x"d4ff4871",
  2038 => x"4f267808",
  2039 => x"48d0ff1e",
  2040 => x"7178e1c8",
  2041 => x"08d4ff48",
  2042 => x"4866c478",
  2043 => x"7808d4ff",
  2044 => x"711e4f26",
  2045 => x"4966c44a",
  2046 => x"ff49721e",
  2047 => x"d0ff87de",
  2048 => x"78e0c048",
  2049 => x"1e4f2626",
  2050 => x"b7c24a71",
  2051 => x"87c303aa",
  2052 => x"ce87c282",
  2053 => x"1e66c482",
  2054 => x"d5ff4972",
  2055 => x"4f262687",
  2056 => x"4ad4ff1e",
  2057 => x"ff7affc3",
  2058 => x"e1c848d0",
  2059 => x"c37ade78",
  2060 => x"7abfd3c5",
  2061 => x"28c84849",
  2062 => x"48717a70",
  2063 => x"7a7028d0",
  2064 => x"28d84871",
  2065 => x"c5c37a70",
  2066 => x"497abfd7",
  2067 => x"7028c848",
  2068 => x"d048717a",
  2069 => x"717a7028",
  2070 => x"7028d848",
  2071 => x"48d0ff7a",
  2072 => x"2678e0c0",
  2073 => x"1e731e4f",
  2074 => x"c5c34a71",
  2075 => x"724bbfd3",
  2076 => x"aae0c02b",
  2077 => x"7287ce04",
  2078 => x"89e0c049",
  2079 => x"bfd7c5c3",
  2080 => x"cf2b714b",
  2081 => x"49e0c087",
  2082 => x"c5c38972",
  2083 => x"7148bfd7",
  2084 => x"b3497030",
  2085 => x"739b66c8",
  2086 => x"2687c448",
  2087 => x"264c264d",
  2088 => x"0e4f264b",
  2089 => x"5d5c5b5e",
  2090 => x"7186ec0e",
  2091 => x"d3c5c34b",
  2092 => x"734c7ebf",
  2093 => x"abe0c02c",
  2094 => x"87e0c004",
  2095 => x"c048a6c4",
  2096 => x"c0497378",
  2097 => x"4a7189e0",
  2098 => x"4866e4c0",
  2099 => x"a6cc3072",
  2100 => x"d7c5c358",
  2101 => x"714c4dbf",
  2102 => x"87e4c02c",
  2103 => x"e4c04973",
  2104 => x"30714866",
  2105 => x"c058a6c8",
  2106 => x"897349e0",
  2107 => x"4866e4c0",
  2108 => x"a6cc2871",
  2109 => x"d7c5c358",
  2110 => x"71484dbf",
  2111 => x"b4497030",
  2112 => x"9c66e4c0",
  2113 => x"e8c084c1",
  2114 => x"c204ac66",
  2115 => x"c04cc087",
  2116 => x"d304abe0",
  2117 => x"48a6cc87",
  2118 => x"497378c0",
  2119 => x"7489e0c0",
  2120 => x"d4307148",
  2121 => x"87d558a6",
  2122 => x"48744973",
  2123 => x"a6d03071",
  2124 => x"49e0c058",
  2125 => x"48748973",
  2126 => x"a6d42871",
  2127 => x"4a66c458",
  2128 => x"9a6ebaff",
  2129 => x"ff4966c8",
  2130 => x"729975b9",
  2131 => x"b066cc48",
  2132 => x"58d7c5c3",
  2133 => x"66d04871",
  2134 => x"dbc5c3b0",
  2135 => x"87c0fb58",
  2136 => x"f6fc8eec",
  2137 => x"d0ff1e87",
  2138 => x"78c9c848",
  2139 => x"d4ff4871",
  2140 => x"4f267808",
  2141 => x"494a711e",
  2142 => x"d0ff87eb",
  2143 => x"2678c848",
  2144 => x"1e731e4f",
  2145 => x"c5c34b71",
  2146 => x"c302bfe7",
  2147 => x"87ebc287",
  2148 => x"c848d0ff",
  2149 => x"497378c9",
  2150 => x"ffb1e0c0",
  2151 => x"787148d4",
  2152 => x"48dbc5c3",
  2153 => x"66c878c0",
  2154 => x"c387c502",
  2155 => x"87c249ff",
  2156 => x"c5c349c0",
  2157 => x"66cc59e3",
  2158 => x"c587c602",
  2159 => x"c44ad5d5",
  2160 => x"ffffcf87",
  2161 => x"e7c5c34a",
  2162 => x"e7c5c35a",
  2163 => x"c478c148",
  2164 => x"264d2687",
  2165 => x"264b264c",
  2166 => x"5b5e0e4f",
  2167 => x"710e5d5c",
  2168 => x"e3c5c34a",
  2169 => x"9a724cbf",
  2170 => x"4987cb02",
  2171 => x"c5c291c8",
  2172 => x"83714bf7",
  2173 => x"c9c287c4",
  2174 => x"4dc04bf7",
  2175 => x"99744913",
  2176 => x"bfdfc5c3",
  2177 => x"48d4ffb9",
  2178 => x"b7c17871",
  2179 => x"b7c8852c",
  2180 => x"87e804ad",
  2181 => x"bfdbc5c3",
  2182 => x"c380c848",
  2183 => x"fe58dfc5",
  2184 => x"731e87ef",
  2185 => x"134b711e",
  2186 => x"cb029a4a",
  2187 => x"fe497287",
  2188 => x"4a1387e7",
  2189 => x"87f5059a",
  2190 => x"1e87dafe",
  2191 => x"bfdbc5c3",
  2192 => x"dbc5c349",
  2193 => x"78a1c148",
  2194 => x"a9b7c0c4",
  2195 => x"ff87db03",
  2196 => x"c5c348d4",
  2197 => x"c378bfdf",
  2198 => x"49bfdbc5",
  2199 => x"48dbc5c3",
  2200 => x"c478a1c1",
  2201 => x"04a9b7c0",
  2202 => x"d0ff87e5",
  2203 => x"c378c848",
  2204 => x"c048e7c5",
  2205 => x"004f2678",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"5f5f0000",
  2209 => x"00000000",
  2210 => x"03000303",
  2211 => x"14000003",
  2212 => x"7f147f7f",
  2213 => x"0000147f",
  2214 => x"6b6b2e24",
  2215 => x"4c00123a",
  2216 => x"6c18366a",
  2217 => x"30003256",
  2218 => x"77594f7e",
  2219 => x"0040683a",
  2220 => x"03070400",
  2221 => x"00000000",
  2222 => x"633e1c00",
  2223 => x"00000041",
  2224 => x"3e634100",
  2225 => x"0800001c",
  2226 => x"1c1c3e2a",
  2227 => x"00082a3e",
  2228 => x"3e3e0808",
  2229 => x"00000808",
  2230 => x"60e08000",
  2231 => x"00000000",
  2232 => x"08080808",
  2233 => x"00000808",
  2234 => x"60600000",
  2235 => x"40000000",
  2236 => x"0c183060",
  2237 => x"00010306",
  2238 => x"4d597f3e",
  2239 => x"00003e7f",
  2240 => x"7f7f0604",
  2241 => x"00000000",
  2242 => x"59716342",
  2243 => x"0000464f",
  2244 => x"49496322",
  2245 => x"1800367f",
  2246 => x"7f13161c",
  2247 => x"0000107f",
  2248 => x"45456727",
  2249 => x"0000397d",
  2250 => x"494b7e3c",
  2251 => x"00003079",
  2252 => x"79710101",
  2253 => x"0000070f",
  2254 => x"49497f36",
  2255 => x"0000367f",
  2256 => x"69494f06",
  2257 => x"00001e3f",
  2258 => x"66660000",
  2259 => x"00000000",
  2260 => x"66e68000",
  2261 => x"00000000",
  2262 => x"14140808",
  2263 => x"00002222",
  2264 => x"14141414",
  2265 => x"00001414",
  2266 => x"14142222",
  2267 => x"00000808",
  2268 => x"59510302",
  2269 => x"3e00060f",
  2270 => x"555d417f",
  2271 => x"00001e1f",
  2272 => x"09097f7e",
  2273 => x"00007e7f",
  2274 => x"49497f7f",
  2275 => x"0000367f",
  2276 => x"41633e1c",
  2277 => x"00004141",
  2278 => x"63417f7f",
  2279 => x"00001c3e",
  2280 => x"49497f7f",
  2281 => x"00004141",
  2282 => x"09097f7f",
  2283 => x"00000101",
  2284 => x"49417f3e",
  2285 => x"00007a7b",
  2286 => x"08087f7f",
  2287 => x"00007f7f",
  2288 => x"7f7f4100",
  2289 => x"00000041",
  2290 => x"40406020",
  2291 => x"7f003f7f",
  2292 => x"361c087f",
  2293 => x"00004163",
  2294 => x"40407f7f",
  2295 => x"7f004040",
  2296 => x"060c067f",
  2297 => x"7f007f7f",
  2298 => x"180c067f",
  2299 => x"00007f7f",
  2300 => x"41417f3e",
  2301 => x"00003e7f",
  2302 => x"09097f7f",
  2303 => x"3e00060f",
  2304 => x"7f61417f",
  2305 => x"0000407e",
  2306 => x"19097f7f",
  2307 => x"0000667f",
  2308 => x"594d6f26",
  2309 => x"0000327b",
  2310 => x"7f7f0101",
  2311 => x"00000101",
  2312 => x"40407f3f",
  2313 => x"00003f7f",
  2314 => x"70703f0f",
  2315 => x"7f000f3f",
  2316 => x"3018307f",
  2317 => x"41007f7f",
  2318 => x"1c1c3663",
  2319 => x"01416336",
  2320 => x"7c7c0603",
  2321 => x"61010306",
  2322 => x"474d5971",
  2323 => x"00004143",
  2324 => x"417f7f00",
  2325 => x"01000041",
  2326 => x"180c0603",
  2327 => x"00406030",
  2328 => x"7f414100",
  2329 => x"0800007f",
  2330 => x"0603060c",
  2331 => x"8000080c",
  2332 => x"80808080",
  2333 => x"00008080",
  2334 => x"07030000",
  2335 => x"00000004",
  2336 => x"54547420",
  2337 => x"0000787c",
  2338 => x"44447f7f",
  2339 => x"0000387c",
  2340 => x"44447c38",
  2341 => x"00000044",
  2342 => x"44447c38",
  2343 => x"00007f7f",
  2344 => x"54547c38",
  2345 => x"0000185c",
  2346 => x"057f7e04",
  2347 => x"00000005",
  2348 => x"a4a4bc18",
  2349 => x"00007cfc",
  2350 => x"04047f7f",
  2351 => x"0000787c",
  2352 => x"7d3d0000",
  2353 => x"00000040",
  2354 => x"fd808080",
  2355 => x"0000007d",
  2356 => x"38107f7f",
  2357 => x"0000446c",
  2358 => x"7f3f0000",
  2359 => x"7c000040",
  2360 => x"0c180c7c",
  2361 => x"0000787c",
  2362 => x"04047c7c",
  2363 => x"0000787c",
  2364 => x"44447c38",
  2365 => x"0000387c",
  2366 => x"2424fcfc",
  2367 => x"0000183c",
  2368 => x"24243c18",
  2369 => x"0000fcfc",
  2370 => x"04047c7c",
  2371 => x"0000080c",
  2372 => x"54545c48",
  2373 => x"00002074",
  2374 => x"447f3f04",
  2375 => x"00000044",
  2376 => x"40407c3c",
  2377 => x"00007c7c",
  2378 => x"60603c1c",
  2379 => x"3c001c3c",
  2380 => x"6030607c",
  2381 => x"44003c7c",
  2382 => x"3810386c",
  2383 => x"0000446c",
  2384 => x"60e0bc1c",
  2385 => x"00001c3c",
  2386 => x"5c746444",
  2387 => x"0000444c",
  2388 => x"773e0808",
  2389 => x"00004141",
  2390 => x"7f7f0000",
  2391 => x"00000000",
  2392 => x"3e774141",
  2393 => x"02000808",
  2394 => x"02030101",
  2395 => x"7f000102",
  2396 => x"7f7f7f7f",
  2397 => x"08007f7f",
  2398 => x"3e1c1c08",
  2399 => x"7f7f7f3e",
  2400 => x"1c3e3e7f",
  2401 => x"0008081c",
  2402 => x"7c7c1810",
  2403 => x"00001018",
  2404 => x"7c7c3010",
  2405 => x"10001030",
  2406 => x"78606030",
  2407 => x"4200061e",
  2408 => x"3c183c66",
  2409 => x"78004266",
  2410 => x"c6c26a38",
  2411 => x"6000386c",
  2412 => x"00600000",
  2413 => x"0e006000",
  2414 => x"5d5c5b5e",
  2415 => x"4c711e0e",
  2416 => x"bff8c5c3",
  2417 => x"c04bc04d",
  2418 => x"02ab741e",
  2419 => x"a6c487c7",
  2420 => x"c578c048",
  2421 => x"48a6c487",
  2422 => x"66c478c1",
  2423 => x"ee49731e",
  2424 => x"86c887df",
  2425 => x"ef49e0c0",
  2426 => x"a5c487ef",
  2427 => x"f0496a4a",
  2428 => x"c6f187f0",
  2429 => x"c185cb87",
  2430 => x"abb7c883",
  2431 => x"87c7ff04",
  2432 => x"264d2626",
  2433 => x"264b264c",
  2434 => x"4a711e4f",
  2435 => x"5afcc5c3",
  2436 => x"48fcc5c3",
  2437 => x"fe4978c7",
  2438 => x"4f2687dd",
  2439 => x"711e731e",
  2440 => x"aab7c04a",
  2441 => x"c287d303",
  2442 => x"05bffbe5",
  2443 => x"4bc187c4",
  2444 => x"4bc087c2",
  2445 => x"5bffe5c2",
  2446 => x"e5c287c4",
  2447 => x"e5c25aff",
  2448 => x"c14abffb",
  2449 => x"a2c0c19a",
  2450 => x"87e8ec49",
  2451 => x"e5c248fc",
  2452 => x"fe78bffb",
  2453 => x"711e87ef",
  2454 => x"1e66c44a",
  2455 => x"e6e64972",
  2456 => x"4f262687",
  2457 => x"fbe5c21e",
  2458 => x"daff49bf",
  2459 => x"c5c387f6",
  2460 => x"bfe848f0",
  2461 => x"ecc5c378",
  2462 => x"78bfec48",
  2463 => x"bff0c5c3",
  2464 => x"ffc3494a",
  2465 => x"2ab7c899",
  2466 => x"b0714872",
  2467 => x"58f8c5c3",
  2468 => x"5e0e4f26",
  2469 => x"0e5d5c5b",
  2470 => x"c7ff4b71",
  2471 => x"ebc5c387",
  2472 => x"7350c048",
  2473 => x"dbdaff49",
  2474 => x"4c497087",
  2475 => x"eecb9cc2",
  2476 => x"87cfcb49",
  2477 => x"c34d4970",
  2478 => x"bf97ebc5",
  2479 => x"87e4c105",
  2480 => x"c34966d0",
  2481 => x"99bff4c5",
  2482 => x"d487d705",
  2483 => x"c5c34966",
  2484 => x"0599bfec",
  2485 => x"497387cc",
  2486 => x"87e8d9ff",
  2487 => x"c1029870",
  2488 => x"4cc187c2",
  2489 => x"7587fdfd",
  2490 => x"87e3ca49",
  2491 => x"c6029870",
  2492 => x"ebc5c387",
  2493 => x"c350c148",
  2494 => x"bf97ebc5",
  2495 => x"87e4c005",
  2496 => x"bff4c5c3",
  2497 => x"9966d049",
  2498 => x"87d6ff05",
  2499 => x"bfecc5c3",
  2500 => x"9966d449",
  2501 => x"87caff05",
  2502 => x"d8ff4973",
  2503 => x"987087e6",
  2504 => x"87fefe05",
  2505 => x"d8fb4874",
  2506 => x"5b5e0e87",
  2507 => x"f40e5d5c",
  2508 => x"4c4dc086",
  2509 => x"c47ebfec",
  2510 => x"c5c348a6",
  2511 => x"c178bff8",
  2512 => x"c71ec01e",
  2513 => x"87cafd49",
  2514 => x"987086c8",
  2515 => x"ff87ce02",
  2516 => x"87c8fb49",
  2517 => x"ff49dac1",
  2518 => x"c187e9d7",
  2519 => x"ebc5c34d",
  2520 => x"c302bf97",
  2521 => x"87ccd587",
  2522 => x"bff0c5c3",
  2523 => x"fbe5c24b",
  2524 => x"ebc005bf",
  2525 => x"49fdc387",
  2526 => x"87c8d7ff",
  2527 => x"ff49fac3",
  2528 => x"7387c1d7",
  2529 => x"99ffc349",
  2530 => x"49c01e71",
  2531 => x"7387c7fb",
  2532 => x"29b7c849",
  2533 => x"49c11e71",
  2534 => x"c887fbfa",
  2535 => x"87c1c686",
  2536 => x"bff4c5c3",
  2537 => x"dd029b4b",
  2538 => x"f7e5c287",
  2539 => x"dec749bf",
  2540 => x"05987087",
  2541 => x"4bc087c4",
  2542 => x"e0c287d2",
  2543 => x"87c3c749",
  2544 => x"58fbe5c2",
  2545 => x"e5c287c6",
  2546 => x"78c048f7",
  2547 => x"99c24973",
  2548 => x"c387ce05",
  2549 => x"d5ff49eb",
  2550 => x"497087ea",
  2551 => x"c20299c2",
  2552 => x"734cfb87",
  2553 => x"0599c149",
  2554 => x"f4c387ce",
  2555 => x"d3d5ff49",
  2556 => x"c2497087",
  2557 => x"87c20299",
  2558 => x"49734cfa",
  2559 => x"ce0599c8",
  2560 => x"49f5c387",
  2561 => x"87fcd4ff",
  2562 => x"99c24970",
  2563 => x"c387d502",
  2564 => x"02bffcc5",
  2565 => x"c14887ca",
  2566 => x"c0c6c388",
  2567 => x"87c2c058",
  2568 => x"4dc14cff",
  2569 => x"99c44973",
  2570 => x"c387ce05",
  2571 => x"d4ff49f2",
  2572 => x"497087d2",
  2573 => x"dc0299c2",
  2574 => x"fcc5c387",
  2575 => x"c7487ebf",
  2576 => x"c003a8b7",
  2577 => x"486e87cb",
  2578 => x"c6c380c1",
  2579 => x"c2c058c0",
  2580 => x"c14cfe87",
  2581 => x"49fdc34d",
  2582 => x"87e8d3ff",
  2583 => x"99c24970",
  2584 => x"87d5c002",
  2585 => x"bffcc5c3",
  2586 => x"87c9c002",
  2587 => x"48fcc5c3",
  2588 => x"c2c078c0",
  2589 => x"c14cfd87",
  2590 => x"49fac34d",
  2591 => x"87c4d3ff",
  2592 => x"99c24970",
  2593 => x"87d9c002",
  2594 => x"bffcc5c3",
  2595 => x"a8b7c748",
  2596 => x"87c9c003",
  2597 => x"48fcc5c3",
  2598 => x"c2c078c7",
  2599 => x"c14cfc87",
  2600 => x"acb7c04d",
  2601 => x"87d1c003",
  2602 => x"c14a66c4",
  2603 => x"026a82d8",
  2604 => x"6a87c6c0",
  2605 => x"7349744b",
  2606 => x"c31ec00f",
  2607 => x"dac11ef0",
  2608 => x"87cef749",
  2609 => x"987086c8",
  2610 => x"87e2c002",
  2611 => x"c348a6c8",
  2612 => x"78bffcc5",
  2613 => x"cb4966c8",
  2614 => x"4866c491",
  2615 => x"7e708071",
  2616 => x"c002bf6e",
  2617 => x"bf6e87c8",
  2618 => x"4966c84b",
  2619 => x"9d750f73",
  2620 => x"87c8c002",
  2621 => x"bffcc5c3",
  2622 => x"87fbf249",
  2623 => x"bfffe5c2",
  2624 => x"87ddc002",
  2625 => x"87c7c249",
  2626 => x"c0029870",
  2627 => x"c5c387d3",
  2628 => x"f249bffc",
  2629 => x"49c087e1",
  2630 => x"c287c1f4",
  2631 => x"c048ffe5",
  2632 => x"f38ef478",
  2633 => x"5e0e87db",
  2634 => x"0e5d5c5b",
  2635 => x"c34c711e",
  2636 => x"49bff8c5",
  2637 => x"4da1cdc1",
  2638 => x"6981d1c1",
  2639 => x"029c747e",
  2640 => x"a5c487cf",
  2641 => x"c37b744b",
  2642 => x"49bff8c5",
  2643 => x"6e87faf2",
  2644 => x"059c747b",
  2645 => x"4bc087c4",
  2646 => x"4bc187c2",
  2647 => x"fbf24973",
  2648 => x"0266d487",
  2649 => x"da4987c7",
  2650 => x"c24a7087",
  2651 => x"c24ac087",
  2652 => x"265ac3e6",
  2653 => x"0087caf2",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"1e000000",
  2657 => x"c8ff4a71",
  2658 => x"a17249bf",
  2659 => x"1e4f2648",
  2660 => x"89bfc8ff",
  2661 => x"c0c0c0fe",
  2662 => x"01a9c0c0",
  2663 => x"4ac087c4",
  2664 => x"4ac187c2",
  2665 => x"4f264872",
  2666 => x"5c5b5e0e",
  2667 => x"4b710e5d",
  2668 => x"d04cd4ff",
  2669 => x"78c04866",
  2670 => x"d8ff49d6",
  2671 => x"ffc387cf",
  2672 => x"c3496c7c",
  2673 => x"4d7199ff",
  2674 => x"99f0c349",
  2675 => x"05a9e0c1",
  2676 => x"ffc387cb",
  2677 => x"c3486c7c",
  2678 => x"0866d098",
  2679 => x"7cffc378",
  2680 => x"c8494a6c",
  2681 => x"7cffc331",
  2682 => x"b2714a6c",
  2683 => x"31c84972",
  2684 => x"6c7cffc3",
  2685 => x"72b2714a",
  2686 => x"c331c849",
  2687 => x"4a6c7cff",
  2688 => x"d0ffb271",
  2689 => x"78e0c048",
  2690 => x"c2029b73",
  2691 => x"757b7287",
  2692 => x"264d2648",
  2693 => x"264b264c",
  2694 => x"4f261e4f",
  2695 => x"5c5b5e0e",
  2696 => x"7686f80e",
  2697 => x"49a6c81e",
  2698 => x"c487fdfd",
  2699 => x"6e4b7086",
  2700 => x"03a8c248",
  2701 => x"7387cac3",
  2702 => x"9af0c34a",
  2703 => x"02aad0c1",
  2704 => x"e0c187c7",
  2705 => x"f8c205aa",
  2706 => x"c8497387",
  2707 => x"87c30299",
  2708 => x"7387c6ff",
  2709 => x"c29cc34c",
  2710 => x"cfc105ac",
  2711 => x"4966c487",
  2712 => x"1e7131c9",
  2713 => x"c04a66c4",
  2714 => x"c6c392f8",
  2715 => x"817249c0",
  2716 => x"87eac0fe",
  2717 => x"1e4966c4",
  2718 => x"ff49e3c0",
  2719 => x"d887f3d5",
  2720 => x"c8d5ff49",
  2721 => x"1ec0c887",
  2722 => x"49caf4c2",
  2723 => x"87cbd9fd",
  2724 => x"c048d0ff",
  2725 => x"f4c278e0",
  2726 => x"66d01eca",
  2727 => x"92f8c04a",
  2728 => x"49c0c6c3",
  2729 => x"fbfd8172",
  2730 => x"86d087f3",
  2731 => x"c105acc1",
  2732 => x"66c487cf",
  2733 => x"7131c949",
  2734 => x"4a66c41e",
  2735 => x"c392f8c0",
  2736 => x"7249c0c6",
  2737 => x"d5fffd81",
  2738 => x"caf4c287",
  2739 => x"4a66c81e",
  2740 => x"c392f8c0",
  2741 => x"7249c0c6",
  2742 => x"fdf9fd81",
  2743 => x"4966c887",
  2744 => x"49e3c01e",
  2745 => x"87cad4ff",
  2746 => x"d3ff49d7",
  2747 => x"c0c887df",
  2748 => x"caf4c21e",
  2749 => x"ccd7fd49",
  2750 => x"ff86d087",
  2751 => x"e0c048d0",
  2752 => x"fc8ef878",
  2753 => x"5e0e87cd",
  2754 => x"0e5d5c5b",
  2755 => x"ff4d711e",
  2756 => x"66d44cd4",
  2757 => x"b7c3487e",
  2758 => x"87c506a8",
  2759 => x"e3c148c0",
  2760 => x"fe497587",
  2761 => x"7587efcf",
  2762 => x"4b66c41e",
  2763 => x"c393f8c0",
  2764 => x"7383c0c6",
  2765 => x"d4f4fd49",
  2766 => x"6b83c887",
  2767 => x"48d0ff4b",
  2768 => x"dd78e1c8",
  2769 => x"c349737c",
  2770 => x"7c7199ff",
  2771 => x"b7c84973",
  2772 => x"99ffc329",
  2773 => x"49737c71",
  2774 => x"c329b7d0",
  2775 => x"7c7199ff",
  2776 => x"b7d84973",
  2777 => x"c07c7129",
  2778 => x"7c7c7c7c",
  2779 => x"7c7c7c7c",
  2780 => x"7c7c7c7c",
  2781 => x"c478e0c0",
  2782 => x"49dc1e66",
  2783 => x"87f2d1ff",
  2784 => x"487386c8",
  2785 => x"87c9fa26",
  2786 => x"5c5b5e0e",
  2787 => x"711e0e5d",
  2788 => x"4bd4ff7e",
  2789 => x"c7c31e6e",
  2790 => x"f2fd49f0",
  2791 => x"86c487ef",
  2792 => x"029d4d70",
  2793 => x"c387c3c3",
  2794 => x"4cbff8c7",
  2795 => x"cdfe496e",
  2796 => x"d0ff87e4",
  2797 => x"78c5c848",
  2798 => x"c07bd6c1",
  2799 => x"c17b154a",
  2800 => x"b7e0c082",
  2801 => x"87f504aa",
  2802 => x"c448d0ff",
  2803 => x"78c5c878",
  2804 => x"c17bd3c1",
  2805 => x"7478c47b",
  2806 => x"fcc1029c",
  2807 => x"caf4c287",
  2808 => x"4dc0c87e",
  2809 => x"acb7c08c",
  2810 => x"c887c603",
  2811 => x"c04da4c0",
  2812 => x"fbc0c34c",
  2813 => x"d049bf97",
  2814 => x"87d20299",
  2815 => x"c7c31ec0",
  2816 => x"f5fd49f0",
  2817 => x"86c487d4",
  2818 => x"c04a4970",
  2819 => x"f4c287ef",
  2820 => x"c7c31eca",
  2821 => x"f5fd49f0",
  2822 => x"86c487c0",
  2823 => x"ff4a4970",
  2824 => x"c5c848d0",
  2825 => x"7bd4c178",
  2826 => x"7bbf976e",
  2827 => x"80c1486e",
  2828 => x"8dc17e70",
  2829 => x"87f0ff05",
  2830 => x"c448d0ff",
  2831 => x"059a7278",
  2832 => x"48c087c5",
  2833 => x"c187e5c0",
  2834 => x"f0c7c31e",
  2835 => x"e8f2fd49",
  2836 => x"7486c487",
  2837 => x"c4fe059c",
  2838 => x"48d0ff87",
  2839 => x"c178c5c8",
  2840 => x"7bc07bd3",
  2841 => x"48c178c4",
  2842 => x"48c087c2",
  2843 => x"264d2626",
  2844 => x"264b264c",
  2845 => x"5b5e0e4f",
  2846 => x"4b710e5c",
  2847 => x"d80266cc",
  2848 => x"f0c04c87",
  2849 => x"87d8028c",
  2850 => x"8ac14a74",
  2851 => x"8a87d102",
  2852 => x"8a87cd02",
  2853 => x"d787c902",
  2854 => x"fb497387",
  2855 => x"87d087ea",
  2856 => x"49c01e74",
  2857 => x"7487dff9",
  2858 => x"f949731e",
  2859 => x"86c887d8",
  2860 => x"0087fcfe",
  2861 => x"ddf3c21e",
  2862 => x"b9c149bf",
  2863 => x"59e1f3c2",
  2864 => x"c348d4ff",
  2865 => x"d0ff78ff",
  2866 => x"78e1c848",
  2867 => x"c148d4ff",
  2868 => x"7131c478",
  2869 => x"48d0ff78",
  2870 => x"2678e0c0",
  2871 => x"0000004f",
  2872 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
