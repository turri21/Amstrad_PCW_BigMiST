
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"78",x"e0",x"c0",x"48"),
     1 => (x"1e",x"4f",x"26",x"26"),
     2 => (x"b7",x"c2",x"4a",x"71"),
     3 => (x"87",x"c3",x"03",x"aa"),
     4 => (x"ce",x"87",x"c2",x"82"),
     5 => (x"1e",x"66",x"c4",x"82"),
     6 => (x"d5",x"ff",x"49",x"72"),
     7 => (x"4f",x"26",x"26",x"87"),
     8 => (x"4a",x"d4",x"ff",x"1e"),
     9 => (x"ff",x"7a",x"ff",x"c3"),
    10 => (x"e1",x"c8",x"48",x"d0"),
    11 => (x"c3",x"7a",x"de",x"78"),
    12 => (x"7a",x"bf",x"d3",x"c5"),
    13 => (x"28",x"c8",x"48",x"49"),
    14 => (x"48",x"71",x"7a",x"70"),
    15 => (x"7a",x"70",x"28",x"d0"),
    16 => (x"28",x"d8",x"48",x"71"),
    17 => (x"c5",x"c3",x"7a",x"70"),
    18 => (x"49",x"7a",x"bf",x"d7"),
    19 => (x"70",x"28",x"c8",x"48"),
    20 => (x"d0",x"48",x"71",x"7a"),
    21 => (x"71",x"7a",x"70",x"28"),
    22 => (x"70",x"28",x"d8",x"48"),
    23 => (x"48",x"d0",x"ff",x"7a"),
    24 => (x"26",x"78",x"e0",x"c0"),
    25 => (x"1e",x"73",x"1e",x"4f"),
    26 => (x"c5",x"c3",x"4a",x"71"),
    27 => (x"72",x"4b",x"bf",x"d3"),
    28 => (x"aa",x"e0",x"c0",x"2b"),
    29 => (x"72",x"87",x"ce",x"04"),
    30 => (x"89",x"e0",x"c0",x"49"),
    31 => (x"bf",x"d7",x"c5",x"c3"),
    32 => (x"cf",x"2b",x"71",x"4b"),
    33 => (x"49",x"e0",x"c0",x"87"),
    34 => (x"c5",x"c3",x"89",x"72"),
    35 => (x"71",x"48",x"bf",x"d7"),
    36 => (x"b3",x"49",x"70",x"30"),
    37 => (x"73",x"9b",x"66",x"c8"),
    38 => (x"26",x"87",x"c4",x"48"),
    39 => (x"26",x"4c",x"26",x"4d"),
    40 => (x"0e",x"4f",x"26",x"4b"),
    41 => (x"5d",x"5c",x"5b",x"5e"),
    42 => (x"71",x"86",x"ec",x"0e"),
    43 => (x"d3",x"c5",x"c3",x"4b"),
    44 => (x"73",x"4c",x"7e",x"bf"),
    45 => (x"ab",x"e0",x"c0",x"2c"),
    46 => (x"87",x"e0",x"c0",x"04"),
    47 => (x"c0",x"48",x"a6",x"c4"),
    48 => (x"c0",x"49",x"73",x"78"),
    49 => (x"4a",x"71",x"89",x"e0"),
    50 => (x"48",x"66",x"e4",x"c0"),
    51 => (x"a6",x"cc",x"30",x"72"),
    52 => (x"d7",x"c5",x"c3",x"58"),
    53 => (x"71",x"4c",x"4d",x"bf"),
    54 => (x"87",x"e4",x"c0",x"2c"),
    55 => (x"e4",x"c0",x"49",x"73"),
    56 => (x"30",x"71",x"48",x"66"),
    57 => (x"c0",x"58",x"a6",x"c8"),
    58 => (x"89",x"73",x"49",x"e0"),
    59 => (x"48",x"66",x"e4",x"c0"),
    60 => (x"a6",x"cc",x"28",x"71"),
    61 => (x"d7",x"c5",x"c3",x"58"),
    62 => (x"71",x"48",x"4d",x"bf"),
    63 => (x"b4",x"49",x"70",x"30"),
    64 => (x"9c",x"66",x"e4",x"c0"),
    65 => (x"e8",x"c0",x"84",x"c1"),
    66 => (x"c2",x"04",x"ac",x"66"),
    67 => (x"c0",x"4c",x"c0",x"87"),
    68 => (x"d3",x"04",x"ab",x"e0"),
    69 => (x"48",x"a6",x"cc",x"87"),
    70 => (x"49",x"73",x"78",x"c0"),
    71 => (x"74",x"89",x"e0",x"c0"),
    72 => (x"d4",x"30",x"71",x"48"),
    73 => (x"87",x"d5",x"58",x"a6"),
    74 => (x"48",x"74",x"49",x"73"),
    75 => (x"a6",x"d0",x"30",x"71"),
    76 => (x"49",x"e0",x"c0",x"58"),
    77 => (x"48",x"74",x"89",x"73"),
    78 => (x"a6",x"d4",x"28",x"71"),
    79 => (x"4a",x"66",x"c4",x"58"),
    80 => (x"9a",x"6e",x"ba",x"ff"),
    81 => (x"ff",x"49",x"66",x"c8"),
    82 => (x"72",x"99",x"75",x"b9"),
    83 => (x"b0",x"66",x"cc",x"48"),
    84 => (x"58",x"d7",x"c5",x"c3"),
    85 => (x"66",x"d0",x"48",x"71"),
    86 => (x"db",x"c5",x"c3",x"b0"),
    87 => (x"87",x"c0",x"fb",x"58"),
    88 => (x"f6",x"fc",x"8e",x"ec"),
    89 => (x"d0",x"ff",x"1e",x"87"),
    90 => (x"78",x"c9",x"c8",x"48"),
    91 => (x"d4",x"ff",x"48",x"71"),
    92 => (x"4f",x"26",x"78",x"08"),
    93 => (x"49",x"4a",x"71",x"1e"),
    94 => (x"d0",x"ff",x"87",x"eb"),
    95 => (x"26",x"78",x"c8",x"48"),
    96 => (x"1e",x"73",x"1e",x"4f"),
    97 => (x"c5",x"c3",x"4b",x"71"),
    98 => (x"c3",x"02",x"bf",x"e7"),
    99 => (x"87",x"eb",x"c2",x"87"),
   100 => (x"c8",x"48",x"d0",x"ff"),
   101 => (x"49",x"73",x"78",x"c9"),
   102 => (x"ff",x"b1",x"e0",x"c0"),
   103 => (x"78",x"71",x"48",x"d4"),
   104 => (x"48",x"db",x"c5",x"c3"),
   105 => (x"66",x"c8",x"78",x"c0"),
   106 => (x"c3",x"87",x"c5",x"02"),
   107 => (x"87",x"c2",x"49",x"ff"),
   108 => (x"c5",x"c3",x"49",x"c0"),
   109 => (x"66",x"cc",x"59",x"e3"),
   110 => (x"c5",x"87",x"c6",x"02"),
   111 => (x"c4",x"4a",x"d5",x"d5"),
   112 => (x"ff",x"ff",x"cf",x"87"),
   113 => (x"e7",x"c5",x"c3",x"4a"),
   114 => (x"e7",x"c5",x"c3",x"5a"),
   115 => (x"c4",x"78",x"c1",x"48"),
   116 => (x"26",x"4d",x"26",x"87"),
   117 => (x"26",x"4b",x"26",x"4c"),
   118 => (x"5b",x"5e",x"0e",x"4f"),
   119 => (x"71",x"0e",x"5d",x"5c"),
   120 => (x"e3",x"c5",x"c3",x"4a"),
   121 => (x"9a",x"72",x"4c",x"bf"),
   122 => (x"49",x"87",x"cb",x"02"),
   123 => (x"c5",x"c2",x"91",x"c8"),
   124 => (x"83",x"71",x"4b",x"f7"),
   125 => (x"c9",x"c2",x"87",x"c4"),
   126 => (x"4d",x"c0",x"4b",x"f7"),
   127 => (x"99",x"74",x"49",x"13"),
   128 => (x"bf",x"df",x"c5",x"c3"),
   129 => (x"48",x"d4",x"ff",x"b9"),
   130 => (x"b7",x"c1",x"78",x"71"),
   131 => (x"b7",x"c8",x"85",x"2c"),
   132 => (x"87",x"e8",x"04",x"ad"),
   133 => (x"bf",x"db",x"c5",x"c3"),
   134 => (x"c3",x"80",x"c8",x"48"),
   135 => (x"fe",x"58",x"df",x"c5"),
   136 => (x"73",x"1e",x"87",x"ef"),
   137 => (x"13",x"4b",x"71",x"1e"),
   138 => (x"cb",x"02",x"9a",x"4a"),
   139 => (x"fe",x"49",x"72",x"87"),
   140 => (x"4a",x"13",x"87",x"e7"),
   141 => (x"87",x"f5",x"05",x"9a"),
   142 => (x"1e",x"87",x"da",x"fe"),
   143 => (x"bf",x"db",x"c5",x"c3"),
   144 => (x"db",x"c5",x"c3",x"49"),
   145 => (x"78",x"a1",x"c1",x"48"),
   146 => (x"a9",x"b7",x"c0",x"c4"),
   147 => (x"ff",x"87",x"db",x"03"),
   148 => (x"c5",x"c3",x"48",x"d4"),
   149 => (x"c3",x"78",x"bf",x"df"),
   150 => (x"49",x"bf",x"db",x"c5"),
   151 => (x"48",x"db",x"c5",x"c3"),
   152 => (x"c4",x"78",x"a1",x"c1"),
   153 => (x"04",x"a9",x"b7",x"c0"),
   154 => (x"d0",x"ff",x"87",x"e5"),
   155 => (x"c3",x"78",x"c8",x"48"),
   156 => (x"c0",x"48",x"e7",x"c5"),
   157 => (x"00",x"4f",x"26",x"78"),
   158 => (x"00",x"00",x"00",x"00"),
   159 => (x"00",x"00",x"00",x"00"),
   160 => (x"5f",x"5f",x"00",x"00"),
   161 => (x"00",x"00",x"00",x"00"),
   162 => (x"03",x"00",x"03",x"03"),
   163 => (x"14",x"00",x"00",x"03"),
   164 => (x"7f",x"14",x"7f",x"7f"),
   165 => (x"00",x"00",x"14",x"7f"),
   166 => (x"6b",x"6b",x"2e",x"24"),
   167 => (x"4c",x"00",x"12",x"3a"),
   168 => (x"6c",x"18",x"36",x"6a"),
   169 => (x"30",x"00",x"32",x"56"),
   170 => (x"77",x"59",x"4f",x"7e"),
   171 => (x"00",x"40",x"68",x"3a"),
   172 => (x"03",x"07",x"04",x"00"),
   173 => (x"00",x"00",x"00",x"00"),
   174 => (x"63",x"3e",x"1c",x"00"),
   175 => (x"00",x"00",x"00",x"41"),
   176 => (x"3e",x"63",x"41",x"00"),
   177 => (x"08",x"00",x"00",x"1c"),
   178 => (x"1c",x"1c",x"3e",x"2a"),
   179 => (x"00",x"08",x"2a",x"3e"),
   180 => (x"3e",x"3e",x"08",x"08"),
   181 => (x"00",x"00",x"08",x"08"),
   182 => (x"60",x"e0",x"80",x"00"),
   183 => (x"00",x"00",x"00",x"00"),
   184 => (x"08",x"08",x"08",x"08"),
   185 => (x"00",x"00",x"08",x"08"),
   186 => (x"60",x"60",x"00",x"00"),
   187 => (x"40",x"00",x"00",x"00"),
   188 => (x"0c",x"18",x"30",x"60"),
   189 => (x"00",x"01",x"03",x"06"),
   190 => (x"4d",x"59",x"7f",x"3e"),
   191 => (x"00",x"00",x"3e",x"7f"),
   192 => (x"7f",x"7f",x"06",x"04"),
   193 => (x"00",x"00",x"00",x"00"),
   194 => (x"59",x"71",x"63",x"42"),
   195 => (x"00",x"00",x"46",x"4f"),
   196 => (x"49",x"49",x"63",x"22"),
   197 => (x"18",x"00",x"36",x"7f"),
   198 => (x"7f",x"13",x"16",x"1c"),
   199 => (x"00",x"00",x"10",x"7f"),
   200 => (x"45",x"45",x"67",x"27"),
   201 => (x"00",x"00",x"39",x"7d"),
   202 => (x"49",x"4b",x"7e",x"3c"),
   203 => (x"00",x"00",x"30",x"79"),
   204 => (x"79",x"71",x"01",x"01"),
   205 => (x"00",x"00",x"07",x"0f"),
   206 => (x"49",x"49",x"7f",x"36"),
   207 => (x"00",x"00",x"36",x"7f"),
   208 => (x"69",x"49",x"4f",x"06"),
   209 => (x"00",x"00",x"1e",x"3f"),
   210 => (x"66",x"66",x"00",x"00"),
   211 => (x"00",x"00",x"00",x"00"),
   212 => (x"66",x"e6",x"80",x"00"),
   213 => (x"00",x"00",x"00",x"00"),
   214 => (x"14",x"14",x"08",x"08"),
   215 => (x"00",x"00",x"22",x"22"),
   216 => (x"14",x"14",x"14",x"14"),
   217 => (x"00",x"00",x"14",x"14"),
   218 => (x"14",x"14",x"22",x"22"),
   219 => (x"00",x"00",x"08",x"08"),
   220 => (x"59",x"51",x"03",x"02"),
   221 => (x"3e",x"00",x"06",x"0f"),
   222 => (x"55",x"5d",x"41",x"7f"),
   223 => (x"00",x"00",x"1e",x"1f"),
   224 => (x"09",x"09",x"7f",x"7e"),
   225 => (x"00",x"00",x"7e",x"7f"),
   226 => (x"49",x"49",x"7f",x"7f"),
   227 => (x"00",x"00",x"36",x"7f"),
   228 => (x"41",x"63",x"3e",x"1c"),
   229 => (x"00",x"00",x"41",x"41"),
   230 => (x"63",x"41",x"7f",x"7f"),
   231 => (x"00",x"00",x"1c",x"3e"),
   232 => (x"49",x"49",x"7f",x"7f"),
   233 => (x"00",x"00",x"41",x"41"),
   234 => (x"09",x"09",x"7f",x"7f"),
   235 => (x"00",x"00",x"01",x"01"),
   236 => (x"49",x"41",x"7f",x"3e"),
   237 => (x"00",x"00",x"7a",x"7b"),
   238 => (x"08",x"08",x"7f",x"7f"),
   239 => (x"00",x"00",x"7f",x"7f"),
   240 => (x"7f",x"7f",x"41",x"00"),
   241 => (x"00",x"00",x"00",x"41"),
   242 => (x"40",x"40",x"60",x"20"),
   243 => (x"7f",x"00",x"3f",x"7f"),
   244 => (x"36",x"1c",x"08",x"7f"),
   245 => (x"00",x"00",x"41",x"63"),
   246 => (x"40",x"40",x"7f",x"7f"),
   247 => (x"7f",x"00",x"40",x"40"),
   248 => (x"06",x"0c",x"06",x"7f"),
   249 => (x"7f",x"00",x"7f",x"7f"),
   250 => (x"18",x"0c",x"06",x"7f"),
   251 => (x"00",x"00",x"7f",x"7f"),
   252 => (x"41",x"41",x"7f",x"3e"),
   253 => (x"00",x"00",x"3e",x"7f"),
   254 => (x"09",x"09",x"7f",x"7f"),
   255 => (x"3e",x"00",x"06",x"0f"),
   256 => (x"7f",x"61",x"41",x"7f"),
   257 => (x"00",x"00",x"40",x"7e"),
   258 => (x"19",x"09",x"7f",x"7f"),
   259 => (x"00",x"00",x"66",x"7f"),
   260 => (x"59",x"4d",x"6f",x"26"),
   261 => (x"00",x"00",x"32",x"7b"),
   262 => (x"7f",x"7f",x"01",x"01"),
   263 => (x"00",x"00",x"01",x"01"),
   264 => (x"40",x"40",x"7f",x"3f"),
   265 => (x"00",x"00",x"3f",x"7f"),
   266 => (x"70",x"70",x"3f",x"0f"),
   267 => (x"7f",x"00",x"0f",x"3f"),
   268 => (x"30",x"18",x"30",x"7f"),
   269 => (x"41",x"00",x"7f",x"7f"),
   270 => (x"1c",x"1c",x"36",x"63"),
   271 => (x"01",x"41",x"63",x"36"),
   272 => (x"7c",x"7c",x"06",x"03"),
   273 => (x"61",x"01",x"03",x"06"),
   274 => (x"47",x"4d",x"59",x"71"),
   275 => (x"00",x"00",x"41",x"43"),
   276 => (x"41",x"7f",x"7f",x"00"),
   277 => (x"01",x"00",x"00",x"41"),
   278 => (x"18",x"0c",x"06",x"03"),
   279 => (x"00",x"40",x"60",x"30"),
   280 => (x"7f",x"41",x"41",x"00"),
   281 => (x"08",x"00",x"00",x"7f"),
   282 => (x"06",x"03",x"06",x"0c"),
   283 => (x"80",x"00",x"08",x"0c"),
   284 => (x"80",x"80",x"80",x"80"),
   285 => (x"00",x"00",x"80",x"80"),
   286 => (x"07",x"03",x"00",x"00"),
   287 => (x"00",x"00",x"00",x"04"),
   288 => (x"54",x"54",x"74",x"20"),
   289 => (x"00",x"00",x"78",x"7c"),
   290 => (x"44",x"44",x"7f",x"7f"),
   291 => (x"00",x"00",x"38",x"7c"),
   292 => (x"44",x"44",x"7c",x"38"),
   293 => (x"00",x"00",x"00",x"44"),
   294 => (x"44",x"44",x"7c",x"38"),
   295 => (x"00",x"00",x"7f",x"7f"),
   296 => (x"54",x"54",x"7c",x"38"),
   297 => (x"00",x"00",x"18",x"5c"),
   298 => (x"05",x"7f",x"7e",x"04"),
   299 => (x"00",x"00",x"00",x"05"),
   300 => (x"a4",x"a4",x"bc",x"18"),
   301 => (x"00",x"00",x"7c",x"fc"),
   302 => (x"04",x"04",x"7f",x"7f"),
   303 => (x"00",x"00",x"78",x"7c"),
   304 => (x"7d",x"3d",x"00",x"00"),
   305 => (x"00",x"00",x"00",x"40"),
   306 => (x"fd",x"80",x"80",x"80"),
   307 => (x"00",x"00",x"00",x"7d"),
   308 => (x"38",x"10",x"7f",x"7f"),
   309 => (x"00",x"00",x"44",x"6c"),
   310 => (x"7f",x"3f",x"00",x"00"),
   311 => (x"7c",x"00",x"00",x"40"),
   312 => (x"0c",x"18",x"0c",x"7c"),
   313 => (x"00",x"00",x"78",x"7c"),
   314 => (x"04",x"04",x"7c",x"7c"),
   315 => (x"00",x"00",x"78",x"7c"),
   316 => (x"44",x"44",x"7c",x"38"),
   317 => (x"00",x"00",x"38",x"7c"),
   318 => (x"24",x"24",x"fc",x"fc"),
   319 => (x"00",x"00",x"18",x"3c"),
   320 => (x"24",x"24",x"3c",x"18"),
   321 => (x"00",x"00",x"fc",x"fc"),
   322 => (x"04",x"04",x"7c",x"7c"),
   323 => (x"00",x"00",x"08",x"0c"),
   324 => (x"54",x"54",x"5c",x"48"),
   325 => (x"00",x"00",x"20",x"74"),
   326 => (x"44",x"7f",x"3f",x"04"),
   327 => (x"00",x"00",x"00",x"44"),
   328 => (x"40",x"40",x"7c",x"3c"),
   329 => (x"00",x"00",x"7c",x"7c"),
   330 => (x"60",x"60",x"3c",x"1c"),
   331 => (x"3c",x"00",x"1c",x"3c"),
   332 => (x"60",x"30",x"60",x"7c"),
   333 => (x"44",x"00",x"3c",x"7c"),
   334 => (x"38",x"10",x"38",x"6c"),
   335 => (x"00",x"00",x"44",x"6c"),
   336 => (x"60",x"e0",x"bc",x"1c"),
   337 => (x"00",x"00",x"1c",x"3c"),
   338 => (x"5c",x"74",x"64",x"44"),
   339 => (x"00",x"00",x"44",x"4c"),
   340 => (x"77",x"3e",x"08",x"08"),
   341 => (x"00",x"00",x"41",x"41"),
   342 => (x"7f",x"7f",x"00",x"00"),
   343 => (x"00",x"00",x"00",x"00"),
   344 => (x"3e",x"77",x"41",x"41"),
   345 => (x"02",x"00",x"08",x"08"),
   346 => (x"02",x"03",x"01",x"01"),
   347 => (x"7f",x"00",x"01",x"02"),
   348 => (x"7f",x"7f",x"7f",x"7f"),
   349 => (x"08",x"00",x"7f",x"7f"),
   350 => (x"3e",x"1c",x"1c",x"08"),
   351 => (x"7f",x"7f",x"7f",x"3e"),
   352 => (x"1c",x"3e",x"3e",x"7f"),
   353 => (x"00",x"08",x"08",x"1c"),
   354 => (x"7c",x"7c",x"18",x"10"),
   355 => (x"00",x"00",x"10",x"18"),
   356 => (x"7c",x"7c",x"30",x"10"),
   357 => (x"10",x"00",x"10",x"30"),
   358 => (x"78",x"60",x"60",x"30"),
   359 => (x"42",x"00",x"06",x"1e"),
   360 => (x"3c",x"18",x"3c",x"66"),
   361 => (x"78",x"00",x"42",x"66"),
   362 => (x"c6",x"c2",x"6a",x"38"),
   363 => (x"60",x"00",x"38",x"6c"),
   364 => (x"00",x"60",x"00",x"00"),
   365 => (x"0e",x"00",x"60",x"00"),
   366 => (x"5d",x"5c",x"5b",x"5e"),
   367 => (x"4c",x"71",x"1e",x"0e"),
   368 => (x"bf",x"f8",x"c5",x"c3"),
   369 => (x"c0",x"4b",x"c0",x"4d"),
   370 => (x"02",x"ab",x"74",x"1e"),
   371 => (x"a6",x"c4",x"87",x"c7"),
   372 => (x"c5",x"78",x"c0",x"48"),
   373 => (x"48",x"a6",x"c4",x"87"),
   374 => (x"66",x"c4",x"78",x"c1"),
   375 => (x"ee",x"49",x"73",x"1e"),
   376 => (x"86",x"c8",x"87",x"df"),
   377 => (x"ef",x"49",x"e0",x"c0"),
   378 => (x"a5",x"c4",x"87",x"ef"),
   379 => (x"f0",x"49",x"6a",x"4a"),
   380 => (x"c6",x"f1",x"87",x"f0"),
   381 => (x"c1",x"85",x"cb",x"87"),
   382 => (x"ab",x"b7",x"c8",x"83"),
   383 => (x"87",x"c7",x"ff",x"04"),
   384 => (x"26",x"4d",x"26",x"26"),
   385 => (x"26",x"4b",x"26",x"4c"),
   386 => (x"4a",x"71",x"1e",x"4f"),
   387 => (x"5a",x"fc",x"c5",x"c3"),
   388 => (x"48",x"fc",x"c5",x"c3"),
   389 => (x"fe",x"49",x"78",x"c7"),
   390 => (x"4f",x"26",x"87",x"dd"),
   391 => (x"71",x"1e",x"73",x"1e"),
   392 => (x"aa",x"b7",x"c0",x"4a"),
   393 => (x"c2",x"87",x"d3",x"03"),
   394 => (x"05",x"bf",x"fb",x"e5"),
   395 => (x"4b",x"c1",x"87",x"c4"),
   396 => (x"4b",x"c0",x"87",x"c2"),
   397 => (x"5b",x"ff",x"e5",x"c2"),
   398 => (x"e5",x"c2",x"87",x"c4"),
   399 => (x"e5",x"c2",x"5a",x"ff"),
   400 => (x"c1",x"4a",x"bf",x"fb"),
   401 => (x"a2",x"c0",x"c1",x"9a"),
   402 => (x"87",x"e8",x"ec",x"49"),
   403 => (x"e5",x"c2",x"48",x"fc"),
   404 => (x"fe",x"78",x"bf",x"fb"),
   405 => (x"71",x"1e",x"87",x"ef"),
   406 => (x"1e",x"66",x"c4",x"4a"),
   407 => (x"e6",x"e6",x"49",x"72"),
   408 => (x"4f",x"26",x"26",x"87"),
   409 => (x"fb",x"e5",x"c2",x"1e"),
   410 => (x"da",x"ff",x"49",x"bf"),
   411 => (x"c5",x"c3",x"87",x"f6"),
   412 => (x"bf",x"e8",x"48",x"f0"),
   413 => (x"ec",x"c5",x"c3",x"78"),
   414 => (x"78",x"bf",x"ec",x"48"),
   415 => (x"bf",x"f0",x"c5",x"c3"),
   416 => (x"ff",x"c3",x"49",x"4a"),
   417 => (x"2a",x"b7",x"c8",x"99"),
   418 => (x"b0",x"71",x"48",x"72"),
   419 => (x"58",x"f8",x"c5",x"c3"),
   420 => (x"5e",x"0e",x"4f",x"26"),
   421 => (x"0e",x"5d",x"5c",x"5b"),
   422 => (x"c7",x"ff",x"4b",x"71"),
   423 => (x"eb",x"c5",x"c3",x"87"),
   424 => (x"73",x"50",x"c0",x"48"),
   425 => (x"db",x"da",x"ff",x"49"),
   426 => (x"4c",x"49",x"70",x"87"),
   427 => (x"ee",x"cb",x"9c",x"c2"),
   428 => (x"87",x"cf",x"cb",x"49"),
   429 => (x"c3",x"4d",x"49",x"70"),
   430 => (x"bf",x"97",x"eb",x"c5"),
   431 => (x"87",x"e4",x"c1",x"05"),
   432 => (x"c3",x"49",x"66",x"d0"),
   433 => (x"99",x"bf",x"f4",x"c5"),
   434 => (x"d4",x"87",x"d7",x"05"),
   435 => (x"c5",x"c3",x"49",x"66"),
   436 => (x"05",x"99",x"bf",x"ec"),
   437 => (x"49",x"73",x"87",x"cc"),
   438 => (x"87",x"e8",x"d9",x"ff"),
   439 => (x"c1",x"02",x"98",x"70"),
   440 => (x"4c",x"c1",x"87",x"c2"),
   441 => (x"75",x"87",x"fd",x"fd"),
   442 => (x"87",x"e3",x"ca",x"49"),
   443 => (x"c6",x"02",x"98",x"70"),
   444 => (x"eb",x"c5",x"c3",x"87"),
   445 => (x"c3",x"50",x"c1",x"48"),
   446 => (x"bf",x"97",x"eb",x"c5"),
   447 => (x"87",x"e4",x"c0",x"05"),
   448 => (x"bf",x"f4",x"c5",x"c3"),
   449 => (x"99",x"66",x"d0",x"49"),
   450 => (x"87",x"d6",x"ff",x"05"),
   451 => (x"bf",x"ec",x"c5",x"c3"),
   452 => (x"99",x"66",x"d4",x"49"),
   453 => (x"87",x"ca",x"ff",x"05"),
   454 => (x"d8",x"ff",x"49",x"73"),
   455 => (x"98",x"70",x"87",x"e6"),
   456 => (x"87",x"fe",x"fe",x"05"),
   457 => (x"d8",x"fb",x"48",x"74"),
   458 => (x"5b",x"5e",x"0e",x"87"),
   459 => (x"f4",x"0e",x"5d",x"5c"),
   460 => (x"4c",x"4d",x"c0",x"86"),
   461 => (x"c4",x"7e",x"bf",x"ec"),
   462 => (x"c5",x"c3",x"48",x"a6"),
   463 => (x"c1",x"78",x"bf",x"f8"),
   464 => (x"c7",x"1e",x"c0",x"1e"),
   465 => (x"87",x"ca",x"fd",x"49"),
   466 => (x"98",x"70",x"86",x"c8"),
   467 => (x"ff",x"87",x"ce",x"02"),
   468 => (x"87",x"c8",x"fb",x"49"),
   469 => (x"ff",x"49",x"da",x"c1"),
   470 => (x"c1",x"87",x"e9",x"d7"),
   471 => (x"eb",x"c5",x"c3",x"4d"),
   472 => (x"c3",x"02",x"bf",x"97"),
   473 => (x"87",x"cc",x"d5",x"87"),
   474 => (x"bf",x"f0",x"c5",x"c3"),
   475 => (x"fb",x"e5",x"c2",x"4b"),
   476 => (x"eb",x"c0",x"05",x"bf"),
   477 => (x"49",x"fd",x"c3",x"87"),
   478 => (x"87",x"c8",x"d7",x"ff"),
   479 => (x"ff",x"49",x"fa",x"c3"),
   480 => (x"73",x"87",x"c1",x"d7"),
   481 => (x"99",x"ff",x"c3",x"49"),
   482 => (x"49",x"c0",x"1e",x"71"),
   483 => (x"73",x"87",x"c7",x"fb"),
   484 => (x"29",x"b7",x"c8",x"49"),
   485 => (x"49",x"c1",x"1e",x"71"),
   486 => (x"c8",x"87",x"fb",x"fa"),
   487 => (x"87",x"c1",x"c6",x"86"),
   488 => (x"bf",x"f4",x"c5",x"c3"),
   489 => (x"dd",x"02",x"9b",x"4b"),
   490 => (x"f7",x"e5",x"c2",x"87"),
   491 => (x"de",x"c7",x"49",x"bf"),
   492 => (x"05",x"98",x"70",x"87"),
   493 => (x"4b",x"c0",x"87",x"c4"),
   494 => (x"e0",x"c2",x"87",x"d2"),
   495 => (x"87",x"c3",x"c7",x"49"),
   496 => (x"58",x"fb",x"e5",x"c2"),
   497 => (x"e5",x"c2",x"87",x"c6"),
   498 => (x"78",x"c0",x"48",x"f7"),
   499 => (x"99",x"c2",x"49",x"73"),
   500 => (x"c3",x"87",x"ce",x"05"),
   501 => (x"d5",x"ff",x"49",x"eb"),
   502 => (x"49",x"70",x"87",x"ea"),
   503 => (x"c2",x"02",x"99",x"c2"),
   504 => (x"73",x"4c",x"fb",x"87"),
   505 => (x"05",x"99",x"c1",x"49"),
   506 => (x"f4",x"c3",x"87",x"ce"),
   507 => (x"d3",x"d5",x"ff",x"49"),
   508 => (x"c2",x"49",x"70",x"87"),
   509 => (x"87",x"c2",x"02",x"99"),
   510 => (x"49",x"73",x"4c",x"fa"),
   511 => (x"ce",x"05",x"99",x"c8"),
   512 => (x"49",x"f5",x"c3",x"87"),
   513 => (x"87",x"fc",x"d4",x"ff"),
   514 => (x"99",x"c2",x"49",x"70"),
   515 => (x"c3",x"87",x"d5",x"02"),
   516 => (x"02",x"bf",x"fc",x"c5"),
   517 => (x"c1",x"48",x"87",x"ca"),
   518 => (x"c0",x"c6",x"c3",x"88"),
   519 => (x"87",x"c2",x"c0",x"58"),
   520 => (x"4d",x"c1",x"4c",x"ff"),
   521 => (x"99",x"c4",x"49",x"73"),
   522 => (x"c3",x"87",x"ce",x"05"),
   523 => (x"d4",x"ff",x"49",x"f2"),
   524 => (x"49",x"70",x"87",x"d2"),
   525 => (x"dc",x"02",x"99",x"c2"),
   526 => (x"fc",x"c5",x"c3",x"87"),
   527 => (x"c7",x"48",x"7e",x"bf"),
   528 => (x"c0",x"03",x"a8",x"b7"),
   529 => (x"48",x"6e",x"87",x"cb"),
   530 => (x"c6",x"c3",x"80",x"c1"),
   531 => (x"c2",x"c0",x"58",x"c0"),
   532 => (x"c1",x"4c",x"fe",x"87"),
   533 => (x"49",x"fd",x"c3",x"4d"),
   534 => (x"87",x"e8",x"d3",x"ff"),
   535 => (x"99",x"c2",x"49",x"70"),
   536 => (x"87",x"d5",x"c0",x"02"),
   537 => (x"bf",x"fc",x"c5",x"c3"),
   538 => (x"87",x"c9",x"c0",x"02"),
   539 => (x"48",x"fc",x"c5",x"c3"),
   540 => (x"c2",x"c0",x"78",x"c0"),
   541 => (x"c1",x"4c",x"fd",x"87"),
   542 => (x"49",x"fa",x"c3",x"4d"),
   543 => (x"87",x"c4",x"d3",x"ff"),
   544 => (x"99",x"c2",x"49",x"70"),
   545 => (x"87",x"d9",x"c0",x"02"),
   546 => (x"bf",x"fc",x"c5",x"c3"),
   547 => (x"a8",x"b7",x"c7",x"48"),
   548 => (x"87",x"c9",x"c0",x"03"),
   549 => (x"48",x"fc",x"c5",x"c3"),
   550 => (x"c2",x"c0",x"78",x"c7"),
   551 => (x"c1",x"4c",x"fc",x"87"),
   552 => (x"ac",x"b7",x"c0",x"4d"),
   553 => (x"87",x"d1",x"c0",x"03"),
   554 => (x"c1",x"4a",x"66",x"c4"),
   555 => (x"02",x"6a",x"82",x"d8"),
   556 => (x"6a",x"87",x"c6",x"c0"),
   557 => (x"73",x"49",x"74",x"4b"),
   558 => (x"c3",x"1e",x"c0",x"0f"),
   559 => (x"da",x"c1",x"1e",x"f0"),
   560 => (x"87",x"ce",x"f7",x"49"),
   561 => (x"98",x"70",x"86",x"c8"),
   562 => (x"87",x"e2",x"c0",x"02"),
   563 => (x"c3",x"48",x"a6",x"c8"),
   564 => (x"78",x"bf",x"fc",x"c5"),
   565 => (x"cb",x"49",x"66",x"c8"),
   566 => (x"48",x"66",x"c4",x"91"),
   567 => (x"7e",x"70",x"80",x"71"),
   568 => (x"c0",x"02",x"bf",x"6e"),
   569 => (x"bf",x"6e",x"87",x"c8"),
   570 => (x"49",x"66",x"c8",x"4b"),
   571 => (x"9d",x"75",x"0f",x"73"),
   572 => (x"87",x"c8",x"c0",x"02"),
   573 => (x"bf",x"fc",x"c5",x"c3"),
   574 => (x"87",x"fb",x"f2",x"49"),
   575 => (x"bf",x"ff",x"e5",x"c2"),
   576 => (x"87",x"dd",x"c0",x"02"),
   577 => (x"87",x"c7",x"c2",x"49"),
   578 => (x"c0",x"02",x"98",x"70"),
   579 => (x"c5",x"c3",x"87",x"d3"),
   580 => (x"f2",x"49",x"bf",x"fc"),
   581 => (x"49",x"c0",x"87",x"e1"),
   582 => (x"c2",x"87",x"c1",x"f4"),
   583 => (x"c0",x"48",x"ff",x"e5"),
   584 => (x"f3",x"8e",x"f4",x"78"),
   585 => (x"5e",x"0e",x"87",x"db"),
   586 => (x"0e",x"5d",x"5c",x"5b"),
   587 => (x"c3",x"4c",x"71",x"1e"),
   588 => (x"49",x"bf",x"f8",x"c5"),
   589 => (x"4d",x"a1",x"cd",x"c1"),
   590 => (x"69",x"81",x"d1",x"c1"),
   591 => (x"02",x"9c",x"74",x"7e"),
   592 => (x"a5",x"c4",x"87",x"cf"),
   593 => (x"c3",x"7b",x"74",x"4b"),
   594 => (x"49",x"bf",x"f8",x"c5"),
   595 => (x"6e",x"87",x"fa",x"f2"),
   596 => (x"05",x"9c",x"74",x"7b"),
   597 => (x"4b",x"c0",x"87",x"c4"),
   598 => (x"4b",x"c1",x"87",x"c2"),
   599 => (x"fb",x"f2",x"49",x"73"),
   600 => (x"02",x"66",x"d4",x"87"),
   601 => (x"da",x"49",x"87",x"c7"),
   602 => (x"c2",x"4a",x"70",x"87"),
   603 => (x"c2",x"4a",x"c0",x"87"),
   604 => (x"26",x"5a",x"c3",x"e6"),
   605 => (x"00",x"87",x"ca",x"f2"),
   606 => (x"00",x"00",x"00",x"00"),
   607 => (x"00",x"00",x"00",x"00"),
   608 => (x"1e",x"00",x"00",x"00"),
   609 => (x"c8",x"ff",x"4a",x"71"),
   610 => (x"a1",x"72",x"49",x"bf"),
   611 => (x"1e",x"4f",x"26",x"48"),
   612 => (x"89",x"bf",x"c8",x"ff"),
   613 => (x"c0",x"c0",x"c0",x"fe"),
   614 => (x"01",x"a9",x"c0",x"c0"),
   615 => (x"4a",x"c0",x"87",x"c4"),
   616 => (x"4a",x"c1",x"87",x"c2"),
   617 => (x"4f",x"26",x"48",x"72"),
   618 => (x"5c",x"5b",x"5e",x"0e"),
   619 => (x"4b",x"71",x"0e",x"5d"),
   620 => (x"d0",x"4c",x"d4",x"ff"),
   621 => (x"78",x"c0",x"48",x"66"),
   622 => (x"d8",x"ff",x"49",x"d6"),
   623 => (x"ff",x"c3",x"87",x"cf"),
   624 => (x"c3",x"49",x"6c",x"7c"),
   625 => (x"4d",x"71",x"99",x"ff"),
   626 => (x"99",x"f0",x"c3",x"49"),
   627 => (x"05",x"a9",x"e0",x"c1"),
   628 => (x"ff",x"c3",x"87",x"cb"),
   629 => (x"c3",x"48",x"6c",x"7c"),
   630 => (x"08",x"66",x"d0",x"98"),
   631 => (x"7c",x"ff",x"c3",x"78"),
   632 => (x"c8",x"49",x"4a",x"6c"),
   633 => (x"7c",x"ff",x"c3",x"31"),
   634 => (x"b2",x"71",x"4a",x"6c"),
   635 => (x"31",x"c8",x"49",x"72"),
   636 => (x"6c",x"7c",x"ff",x"c3"),
   637 => (x"72",x"b2",x"71",x"4a"),
   638 => (x"c3",x"31",x"c8",x"49"),
   639 => (x"4a",x"6c",x"7c",x"ff"),
   640 => (x"d0",x"ff",x"b2",x"71"),
   641 => (x"78",x"e0",x"c0",x"48"),
   642 => (x"c2",x"02",x"9b",x"73"),
   643 => (x"75",x"7b",x"72",x"87"),
   644 => (x"26",x"4d",x"26",x"48"),
   645 => (x"26",x"4b",x"26",x"4c"),
   646 => (x"4f",x"26",x"1e",x"4f"),
   647 => (x"5c",x"5b",x"5e",x"0e"),
   648 => (x"76",x"86",x"f8",x"0e"),
   649 => (x"49",x"a6",x"c8",x"1e"),
   650 => (x"c4",x"87",x"fd",x"fd"),
   651 => (x"6e",x"4b",x"70",x"86"),
   652 => (x"03",x"a8",x"c2",x"48"),
   653 => (x"73",x"87",x"ca",x"c3"),
   654 => (x"9a",x"f0",x"c3",x"4a"),
   655 => (x"02",x"aa",x"d0",x"c1"),
   656 => (x"e0",x"c1",x"87",x"c7"),
   657 => (x"f8",x"c2",x"05",x"aa"),
   658 => (x"c8",x"49",x"73",x"87"),
   659 => (x"87",x"c3",x"02",x"99"),
   660 => (x"73",x"87",x"c6",x"ff"),
   661 => (x"c2",x"9c",x"c3",x"4c"),
   662 => (x"cf",x"c1",x"05",x"ac"),
   663 => (x"49",x"66",x"c4",x"87"),
   664 => (x"1e",x"71",x"31",x"c9"),
   665 => (x"c0",x"4a",x"66",x"c4"),
   666 => (x"c6",x"c3",x"92",x"f8"),
   667 => (x"81",x"72",x"49",x"c0"),
   668 => (x"87",x"ea",x"c0",x"fe"),
   669 => (x"1e",x"49",x"66",x"c4"),
   670 => (x"ff",x"49",x"e3",x"c0"),
   671 => (x"d8",x"87",x"f3",x"d5"),
   672 => (x"c8",x"d5",x"ff",x"49"),
   673 => (x"1e",x"c0",x"c8",x"87"),
   674 => (x"49",x"ca",x"f4",x"c2"),
   675 => (x"87",x"cb",x"d9",x"fd"),
   676 => (x"c0",x"48",x"d0",x"ff"),
   677 => (x"f4",x"c2",x"78",x"e0"),
   678 => (x"66",x"d0",x"1e",x"ca"),
   679 => (x"92",x"f8",x"c0",x"4a"),
   680 => (x"49",x"c0",x"c6",x"c3"),
   681 => (x"fb",x"fd",x"81",x"72"),
   682 => (x"86",x"d0",x"87",x"f3"),
   683 => (x"c1",x"05",x"ac",x"c1"),
   684 => (x"66",x"c4",x"87",x"cf"),
   685 => (x"71",x"31",x"c9",x"49"),
   686 => (x"4a",x"66",x"c4",x"1e"),
   687 => (x"c3",x"92",x"f8",x"c0"),
   688 => (x"72",x"49",x"c0",x"c6"),
   689 => (x"d5",x"ff",x"fd",x"81"),
   690 => (x"ca",x"f4",x"c2",x"87"),
   691 => (x"4a",x"66",x"c8",x"1e"),
   692 => (x"c3",x"92",x"f8",x"c0"),
   693 => (x"72",x"49",x"c0",x"c6"),
   694 => (x"fd",x"f9",x"fd",x"81"),
   695 => (x"49",x"66",x"c8",x"87"),
   696 => (x"49",x"e3",x"c0",x"1e"),
   697 => (x"87",x"ca",x"d4",x"ff"),
   698 => (x"d3",x"ff",x"49",x"d7"),
   699 => (x"c0",x"c8",x"87",x"df"),
   700 => (x"ca",x"f4",x"c2",x"1e"),
   701 => (x"cc",x"d7",x"fd",x"49"),
   702 => (x"ff",x"86",x"d0",x"87"),
   703 => (x"e0",x"c0",x"48",x"d0"),
   704 => (x"fc",x"8e",x"f8",x"78"),
   705 => (x"5e",x"0e",x"87",x"cd"),
   706 => (x"0e",x"5d",x"5c",x"5b"),
   707 => (x"ff",x"4d",x"71",x"1e"),
   708 => (x"66",x"d4",x"4c",x"d4"),
   709 => (x"b7",x"c3",x"48",x"7e"),
   710 => (x"87",x"c5",x"06",x"a8"),
   711 => (x"e3",x"c1",x"48",x"c0"),
   712 => (x"fe",x"49",x"75",x"87"),
   713 => (x"75",x"87",x"ef",x"cf"),
   714 => (x"4b",x"66",x"c4",x"1e"),
   715 => (x"c3",x"93",x"f8",x"c0"),
   716 => (x"73",x"83",x"c0",x"c6"),
   717 => (x"d4",x"f4",x"fd",x"49"),
   718 => (x"6b",x"83",x"c8",x"87"),
   719 => (x"48",x"d0",x"ff",x"4b"),
   720 => (x"dd",x"78",x"e1",x"c8"),
   721 => (x"c3",x"49",x"73",x"7c"),
   722 => (x"7c",x"71",x"99",x"ff"),
   723 => (x"b7",x"c8",x"49",x"73"),
   724 => (x"99",x"ff",x"c3",x"29"),
   725 => (x"49",x"73",x"7c",x"71"),
   726 => (x"c3",x"29",x"b7",x"d0"),
   727 => (x"7c",x"71",x"99",x"ff"),
   728 => (x"b7",x"d8",x"49",x"73"),
   729 => (x"c0",x"7c",x"71",x"29"),
   730 => (x"7c",x"7c",x"7c",x"7c"),
   731 => (x"7c",x"7c",x"7c",x"7c"),
   732 => (x"7c",x"7c",x"7c",x"7c"),
   733 => (x"c4",x"78",x"e0",x"c0"),
   734 => (x"49",x"dc",x"1e",x"66"),
   735 => (x"87",x"f2",x"d1",x"ff"),
   736 => (x"48",x"73",x"86",x"c8"),
   737 => (x"87",x"c9",x"fa",x"26"),
   738 => (x"5c",x"5b",x"5e",x"0e"),
   739 => (x"71",x"1e",x"0e",x"5d"),
   740 => (x"4b",x"d4",x"ff",x"7e"),
   741 => (x"c7",x"c3",x"1e",x"6e"),
   742 => (x"f2",x"fd",x"49",x"f0"),
   743 => (x"86",x"c4",x"87",x"ef"),
   744 => (x"02",x"9d",x"4d",x"70"),
   745 => (x"c3",x"87",x"c3",x"c3"),
   746 => (x"4c",x"bf",x"f8",x"c7"),
   747 => (x"cd",x"fe",x"49",x"6e"),
   748 => (x"d0",x"ff",x"87",x"e4"),
   749 => (x"78",x"c5",x"c8",x"48"),
   750 => (x"c0",x"7b",x"d6",x"c1"),
   751 => (x"c1",x"7b",x"15",x"4a"),
   752 => (x"b7",x"e0",x"c0",x"82"),
   753 => (x"87",x"f5",x"04",x"aa"),
   754 => (x"c4",x"48",x"d0",x"ff"),
   755 => (x"78",x"c5",x"c8",x"78"),
   756 => (x"c1",x"7b",x"d3",x"c1"),
   757 => (x"74",x"78",x"c4",x"7b"),
   758 => (x"fc",x"c1",x"02",x"9c"),
   759 => (x"ca",x"f4",x"c2",x"87"),
   760 => (x"4d",x"c0",x"c8",x"7e"),
   761 => (x"ac",x"b7",x"c0",x"8c"),
   762 => (x"c8",x"87",x"c6",x"03"),
   763 => (x"c0",x"4d",x"a4",x"c0"),
   764 => (x"fb",x"c0",x"c3",x"4c"),
   765 => (x"d0",x"49",x"bf",x"97"),
   766 => (x"87",x"d2",x"02",x"99"),
   767 => (x"c7",x"c3",x"1e",x"c0"),
   768 => (x"f5",x"fd",x"49",x"f0"),
   769 => (x"86",x"c4",x"87",x"d4"),
   770 => (x"c0",x"4a",x"49",x"70"),
   771 => (x"f4",x"c2",x"87",x"ef"),
   772 => (x"c7",x"c3",x"1e",x"ca"),
   773 => (x"f5",x"fd",x"49",x"f0"),
   774 => (x"86",x"c4",x"87",x"c0"),
   775 => (x"ff",x"4a",x"49",x"70"),
   776 => (x"c5",x"c8",x"48",x"d0"),
   777 => (x"7b",x"d4",x"c1",x"78"),
   778 => (x"7b",x"bf",x"97",x"6e"),
   779 => (x"80",x"c1",x"48",x"6e"),
   780 => (x"8d",x"c1",x"7e",x"70"),
   781 => (x"87",x"f0",x"ff",x"05"),
   782 => (x"c4",x"48",x"d0",x"ff"),
   783 => (x"05",x"9a",x"72",x"78"),
   784 => (x"48",x"c0",x"87",x"c5"),
   785 => (x"c1",x"87",x"e5",x"c0"),
   786 => (x"f0",x"c7",x"c3",x"1e"),
   787 => (x"e8",x"f2",x"fd",x"49"),
   788 => (x"74",x"86",x"c4",x"87"),
   789 => (x"c4",x"fe",x"05",x"9c"),
   790 => (x"48",x"d0",x"ff",x"87"),
   791 => (x"c1",x"78",x"c5",x"c8"),
   792 => (x"7b",x"c0",x"7b",x"d3"),
   793 => (x"48",x"c1",x"78",x"c4"),
   794 => (x"48",x"c0",x"87",x"c2"),
   795 => (x"26",x"4d",x"26",x"26"),
   796 => (x"26",x"4b",x"26",x"4c"),
   797 => (x"5b",x"5e",x"0e",x"4f"),
   798 => (x"4b",x"71",x"0e",x"5c"),
   799 => (x"d8",x"02",x"66",x"cc"),
   800 => (x"f0",x"c0",x"4c",x"87"),
   801 => (x"87",x"d8",x"02",x"8c"),
   802 => (x"8a",x"c1",x"4a",x"74"),
   803 => (x"8a",x"87",x"d1",x"02"),
   804 => (x"8a",x"87",x"cd",x"02"),
   805 => (x"d7",x"87",x"c9",x"02"),
   806 => (x"fb",x"49",x"73",x"87"),
   807 => (x"87",x"d0",x"87",x"ea"),
   808 => (x"49",x"c0",x"1e",x"74"),
   809 => (x"74",x"87",x"df",x"f9"),
   810 => (x"f9",x"49",x"73",x"1e"),
   811 => (x"86",x"c8",x"87",x"d8"),
   812 => (x"00",x"87",x"fc",x"fe"),
   813 => (x"dd",x"f3",x"c2",x"1e"),
   814 => (x"b9",x"c1",x"49",x"bf"),
   815 => (x"59",x"e1",x"f3",x"c2"),
   816 => (x"c3",x"48",x"d4",x"ff"),
   817 => (x"d0",x"ff",x"78",x"ff"),
   818 => (x"78",x"e1",x"c8",x"48"),
   819 => (x"c1",x"48",x"d4",x"ff"),
   820 => (x"71",x"31",x"c4",x"78"),
   821 => (x"48",x"d0",x"ff",x"78"),
   822 => (x"26",x"78",x"e0",x"c0"),
   823 => (x"00",x"00",x"00",x"4f"),
   824 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

